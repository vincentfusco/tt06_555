magic
tech sky130A
magscale 1 2
timestamp 1711057506
<< pwell >>
rect 20908 2162 22408 3520
<< psubdiff >>
rect 20944 3450 21040 3484
rect 22276 3450 22372 3484
rect 20944 3388 20978 3450
rect 22338 3388 22372 3450
rect 20944 2232 20978 2300
rect 22338 2232 22372 2300
rect 20944 2198 21040 2232
rect 22276 2198 22372 2232
<< psubdiffcont >>
rect 21040 3450 22276 3484
rect 20944 2300 20978 3388
rect 22338 2300 22372 3388
rect 21040 2198 22276 2232
<< poly >>
rect 22188 3295 22268 3311
rect 22188 3257 22221 3295
rect 22255 3257 22268 3295
rect 22188 3241 22268 3257
rect 21058 3167 21138 3183
rect 21058 3129 21071 3167
rect 21105 3129 21138 3167
rect 21058 3113 21138 3129
rect 21137 2985 21138 3055
rect 22188 3039 22268 3055
rect 22188 3001 22221 3039
rect 22255 3001 22268 3039
rect 22188 2985 22268 3001
rect 21058 2911 21138 2927
rect 21058 2873 21071 2911
rect 21105 2873 21138 2911
rect 21058 2857 21138 2873
rect 21137 2729 21138 2799
rect 22188 2783 22267 2799
rect 22188 2745 22220 2783
rect 22254 2745 22267 2783
rect 22188 2729 22267 2745
rect 21059 2655 21138 2671
rect 21059 2617 21072 2655
rect 21106 2617 21138 2655
rect 21059 2601 21138 2617
rect 21137 2473 21138 2543
rect 22188 2527 22267 2543
rect 22188 2489 22220 2527
rect 22254 2489 22267 2527
rect 22188 2473 22267 2489
rect 21059 2399 21138 2415
rect 21059 2361 21072 2399
rect 21106 2361 21138 2399
rect 21059 2345 21138 2361
<< polycont >>
rect 22221 3257 22255 3295
rect 21071 3129 21105 3167
rect 22221 3001 22255 3039
rect 21071 2873 21105 2911
rect 22220 2745 22254 2783
rect 21072 2617 21106 2655
rect 22220 2489 22254 2527
rect 21072 2361 21106 2399
<< locali >>
rect 20944 3450 21040 3484
rect 22276 3450 22372 3484
rect 20944 3388 20978 3450
rect 22338 3388 22372 3450
rect 22221 3295 22255 3311
rect 22221 3241 22255 3257
rect 21071 3167 21105 3183
rect 21071 3113 21105 3129
rect 22221 3039 22255 3055
rect 22221 2985 22255 3001
rect 21071 2911 21105 2927
rect 21071 2857 21105 2873
rect 22220 2783 22254 2799
rect 22220 2729 22254 2745
rect 21072 2655 21106 2671
rect 21072 2601 21106 2617
rect 22220 2527 22254 2543
rect 22220 2473 22254 2489
rect 21072 2399 21106 2415
rect 21072 2345 21106 2361
rect 20944 2234 20978 2300
rect 22338 2234 22372 2300
rect 20944 2232 22372 2234
rect 20944 2198 21040 2232
rect 22276 2198 22372 2232
rect 20944 2102 22372 2198
<< viali >>
rect 22221 3257 22255 3295
rect 21071 3129 21105 3167
rect 22221 3001 22255 3039
rect 21071 2873 21105 2911
rect 22220 2745 22254 2783
rect 21072 2617 21106 2655
rect 22220 2489 22254 2527
rect 21072 2361 21106 2399
<< metal1 >>
rect 18500 4218 18700 4418
rect 18500 3818 18700 4018
rect 18500 3418 18700 3618
rect 22214 3295 22270 3392
rect 18500 3018 18700 3218
rect 21056 3167 21112 3264
rect 21056 3129 21071 3167
rect 21105 3129 21112 3167
rect 21056 2911 21112 3129
rect 21056 2873 21071 2911
rect 21105 2873 21112 2911
rect 18500 2618 18700 2818
rect 21056 2655 21112 2873
rect 21056 2617 21072 2655
rect 21106 2617 21112 2655
rect 18500 2218 18700 2418
rect 21056 2399 21112 2617
rect 22214 3257 22221 3295
rect 22255 3257 22270 3295
rect 22214 3039 22270 3257
rect 22214 3001 22221 3039
rect 22255 3001 22270 3039
rect 22214 2783 22270 3001
rect 22214 2745 22220 2783
rect 22254 2745 22270 2783
rect 22214 2527 22270 2745
rect 22214 2489 22220 2527
rect 22254 2489 22270 2527
rect 22214 2472 22270 2489
rect 21056 2361 21072 2399
rect 21106 2361 21112 2399
rect 21056 2344 21112 2361
use sky130_fd_pr__nfet_01v8_lvt_Q8GSR7  sky130_fd_pr__nfet_01v8_lvt_Q8GSR7_0
timestamp 1711041017
transform 0 1 21663 -1 0 3084
box -285 -526 285 526
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_diode_left
timestamp 1711041810
transform 0 1 20248 -1 0 1874
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_Q8GSR7  XMn_inp
timestamp 1711041017
transform 0 1 21663 -1 0 2572
box -285 -526 285 526
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_out
timestamp 1711041810
transform 0 1 23036 -1 0 1874
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_tail
timestamp 1711041810
transform 0 1 21642 -1 0 1874
box -296 -734 296 766
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_cs_left
timestamp 1711036998
transform 0 1 20492 -1 0 4456
box -296 -1219 296 1219
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_cs_right
timestamp 1711036998
transform 0 1 22824 -1 0 4456
box -296 -1219 296 1219
use sky130_fd_pr__pfet_01v8_lvt_5VNMZ8  XMp_diode_left
timestamp 1711036998
transform 0 1 20692 -1 0 3866
box -296 -1019 296 1019
use sky130_fd_pr__pfet_01v8_lvt_5VNMZ8  XMp_diode_right
timestamp 1711036998
transform 0 1 22624 -1 0 3866
box -296 -1019 296 1019
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_out_left_top
timestamp 1711036998
transform 0 -1 20492 1 0 4942
box -296 -1219 296 1219
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_out_right_top
timestamp 1711036998
transform 0 -1 22824 1 0 4942
box -296 -1219 296 1219
<< labels >>
flabel metal1 18500 4218 18700 4418 0 FreeSans 256 0 0 0 INp
port 0 nsew
flabel metal1 18500 3818 18700 4018 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 18500 2618 18700 2818 0 FreeSans 256 0 0 0 INn
port 4 nsew
flabel metal1 18500 2218 18700 2418 0 FreeSans 256 0 0 0 bias_n
port 5 nsew
flabel metal1 18500 4218 18700 4418 0 FreeSans 256 0 0 0 vinp
flabel metal1 18500 3818 18700 4018 0 FreeSans 256 0 0 0 vout
flabel metal1 18500 3418 18700 3618 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 18500 3018 18700 3218 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 18500 2618 18700 2818 0 FreeSans 256 0 0 0 vinn
flabel metal1 18500 2218 18700 2418 0 FreeSans 256 0 0 0 vbias_n
<< end >>
