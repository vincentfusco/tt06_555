magic
tech sky130A
magscale 1 2
timestamp 1710860902
<< error_p >>
rect -173 2835 -115 2841
rect 19 2835 77 2841
rect -173 2801 -161 2835
rect 19 2801 31 2835
rect -173 2795 -115 2801
rect 19 2795 77 2801
rect -77 2225 -19 2231
rect 115 2225 173 2231
rect -77 2191 -65 2225
rect 115 2191 127 2225
rect -77 2185 -19 2191
rect 115 2185 173 2191
rect -77 2117 -19 2123
rect 115 2117 173 2123
rect -77 2083 -65 2117
rect 115 2083 127 2117
rect -77 2077 -19 2083
rect 115 2077 173 2083
rect -173 1507 -115 1513
rect 19 1507 77 1513
rect -173 1473 -161 1507
rect 19 1473 31 1507
rect -173 1467 -115 1473
rect 19 1467 77 1473
rect -173 1399 -115 1405
rect 19 1399 77 1405
rect -173 1365 -161 1399
rect 19 1365 31 1399
rect -173 1359 -115 1365
rect 19 1359 77 1365
rect -77 789 -19 795
rect 115 789 173 795
rect -77 755 -65 789
rect 115 755 127 789
rect -77 749 -19 755
rect 115 749 173 755
rect -77 681 -19 687
rect 115 681 173 687
rect -77 647 -65 681
rect 115 647 127 681
rect -77 641 -19 647
rect 115 641 173 647
rect -173 71 -115 77
rect 19 71 77 77
rect -173 37 -161 71
rect 19 37 31 71
rect -173 31 -115 37
rect 19 31 77 37
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect -77 -647 -19 -641
rect 115 -647 173 -641
rect -77 -681 -65 -647
rect 115 -681 127 -647
rect -77 -687 -19 -681
rect 115 -687 173 -681
rect -77 -755 -19 -749
rect 115 -755 173 -749
rect -77 -789 -65 -755
rect 115 -789 127 -755
rect -77 -795 -19 -789
rect 115 -795 173 -789
rect -173 -1365 -115 -1359
rect 19 -1365 77 -1359
rect -173 -1399 -161 -1365
rect 19 -1399 31 -1365
rect -173 -1405 -115 -1399
rect 19 -1405 77 -1399
rect -173 -1473 -115 -1467
rect 19 -1473 77 -1467
rect -173 -1507 -161 -1473
rect 19 -1507 31 -1473
rect -173 -1513 -115 -1507
rect 19 -1513 77 -1507
rect -77 -2083 -19 -2077
rect 115 -2083 173 -2077
rect -77 -2117 -65 -2083
rect 115 -2117 127 -2083
rect -77 -2123 -19 -2117
rect 115 -2123 173 -2117
rect -77 -2191 -19 -2185
rect 115 -2191 173 -2185
rect -77 -2225 -65 -2191
rect 115 -2225 127 -2191
rect -77 -2231 -19 -2225
rect 115 -2231 173 -2225
rect -173 -2801 -115 -2795
rect 19 -2801 77 -2795
rect -173 -2835 -161 -2801
rect 19 -2835 31 -2801
rect -173 -2841 -115 -2835
rect 19 -2841 77 -2835
<< pwell >>
rect -359 -2973 359 2973
<< nmos >>
rect -159 2263 -129 2763
rect -63 2263 -33 2763
rect 33 2263 63 2763
rect 129 2263 159 2763
rect -159 1545 -129 2045
rect -63 1545 -33 2045
rect 33 1545 63 2045
rect 129 1545 159 2045
rect -159 827 -129 1327
rect -63 827 -33 1327
rect 33 827 63 1327
rect 129 827 159 1327
rect -159 109 -129 609
rect -63 109 -33 609
rect 33 109 63 609
rect 129 109 159 609
rect -159 -609 -129 -109
rect -63 -609 -33 -109
rect 33 -609 63 -109
rect 129 -609 159 -109
rect -159 -1327 -129 -827
rect -63 -1327 -33 -827
rect 33 -1327 63 -827
rect 129 -1327 159 -827
rect -159 -2045 -129 -1545
rect -63 -2045 -33 -1545
rect 33 -2045 63 -1545
rect 129 -2045 159 -1545
rect -159 -2763 -129 -2263
rect -63 -2763 -33 -2263
rect 33 -2763 63 -2263
rect 129 -2763 159 -2263
<< ndiff >>
rect -221 2751 -159 2763
rect -221 2275 -209 2751
rect -175 2275 -159 2751
rect -221 2263 -159 2275
rect -129 2751 -63 2763
rect -129 2275 -113 2751
rect -79 2275 -63 2751
rect -129 2263 -63 2275
rect -33 2751 33 2763
rect -33 2275 -17 2751
rect 17 2275 33 2751
rect -33 2263 33 2275
rect 63 2751 129 2763
rect 63 2275 79 2751
rect 113 2275 129 2751
rect 63 2263 129 2275
rect 159 2751 221 2763
rect 159 2275 175 2751
rect 209 2275 221 2751
rect 159 2263 221 2275
rect -221 2033 -159 2045
rect -221 1557 -209 2033
rect -175 1557 -159 2033
rect -221 1545 -159 1557
rect -129 2033 -63 2045
rect -129 1557 -113 2033
rect -79 1557 -63 2033
rect -129 1545 -63 1557
rect -33 2033 33 2045
rect -33 1557 -17 2033
rect 17 1557 33 2033
rect -33 1545 33 1557
rect 63 2033 129 2045
rect 63 1557 79 2033
rect 113 1557 129 2033
rect 63 1545 129 1557
rect 159 2033 221 2045
rect 159 1557 175 2033
rect 209 1557 221 2033
rect 159 1545 221 1557
rect -221 1315 -159 1327
rect -221 839 -209 1315
rect -175 839 -159 1315
rect -221 827 -159 839
rect -129 1315 -63 1327
rect -129 839 -113 1315
rect -79 839 -63 1315
rect -129 827 -63 839
rect -33 1315 33 1327
rect -33 839 -17 1315
rect 17 839 33 1315
rect -33 827 33 839
rect 63 1315 129 1327
rect 63 839 79 1315
rect 113 839 129 1315
rect 63 827 129 839
rect 159 1315 221 1327
rect 159 839 175 1315
rect 209 839 221 1315
rect 159 827 221 839
rect -221 597 -159 609
rect -221 121 -209 597
rect -175 121 -159 597
rect -221 109 -159 121
rect -129 597 -63 609
rect -129 121 -113 597
rect -79 121 -63 597
rect -129 109 -63 121
rect -33 597 33 609
rect -33 121 -17 597
rect 17 121 33 597
rect -33 109 33 121
rect 63 597 129 609
rect 63 121 79 597
rect 113 121 129 597
rect 63 109 129 121
rect 159 597 221 609
rect 159 121 175 597
rect 209 121 221 597
rect 159 109 221 121
rect -221 -121 -159 -109
rect -221 -597 -209 -121
rect -175 -597 -159 -121
rect -221 -609 -159 -597
rect -129 -121 -63 -109
rect -129 -597 -113 -121
rect -79 -597 -63 -121
rect -129 -609 -63 -597
rect -33 -121 33 -109
rect -33 -597 -17 -121
rect 17 -597 33 -121
rect -33 -609 33 -597
rect 63 -121 129 -109
rect 63 -597 79 -121
rect 113 -597 129 -121
rect 63 -609 129 -597
rect 159 -121 221 -109
rect 159 -597 175 -121
rect 209 -597 221 -121
rect 159 -609 221 -597
rect -221 -839 -159 -827
rect -221 -1315 -209 -839
rect -175 -1315 -159 -839
rect -221 -1327 -159 -1315
rect -129 -839 -63 -827
rect -129 -1315 -113 -839
rect -79 -1315 -63 -839
rect -129 -1327 -63 -1315
rect -33 -839 33 -827
rect -33 -1315 -17 -839
rect 17 -1315 33 -839
rect -33 -1327 33 -1315
rect 63 -839 129 -827
rect 63 -1315 79 -839
rect 113 -1315 129 -839
rect 63 -1327 129 -1315
rect 159 -839 221 -827
rect 159 -1315 175 -839
rect 209 -1315 221 -839
rect 159 -1327 221 -1315
rect -221 -1557 -159 -1545
rect -221 -2033 -209 -1557
rect -175 -2033 -159 -1557
rect -221 -2045 -159 -2033
rect -129 -1557 -63 -1545
rect -129 -2033 -113 -1557
rect -79 -2033 -63 -1557
rect -129 -2045 -63 -2033
rect -33 -1557 33 -1545
rect -33 -2033 -17 -1557
rect 17 -2033 33 -1557
rect -33 -2045 33 -2033
rect 63 -1557 129 -1545
rect 63 -2033 79 -1557
rect 113 -2033 129 -1557
rect 63 -2045 129 -2033
rect 159 -1557 221 -1545
rect 159 -2033 175 -1557
rect 209 -2033 221 -1557
rect 159 -2045 221 -2033
rect -221 -2275 -159 -2263
rect -221 -2751 -209 -2275
rect -175 -2751 -159 -2275
rect -221 -2763 -159 -2751
rect -129 -2275 -63 -2263
rect -129 -2751 -113 -2275
rect -79 -2751 -63 -2275
rect -129 -2763 -63 -2751
rect -33 -2275 33 -2263
rect -33 -2751 -17 -2275
rect 17 -2751 33 -2275
rect -33 -2763 33 -2751
rect 63 -2275 129 -2263
rect 63 -2751 79 -2275
rect 113 -2751 129 -2275
rect 63 -2763 129 -2751
rect 159 -2275 221 -2263
rect 159 -2751 175 -2275
rect 209 -2751 221 -2275
rect 159 -2763 221 -2751
<< ndiffc >>
rect -209 2275 -175 2751
rect -113 2275 -79 2751
rect -17 2275 17 2751
rect 79 2275 113 2751
rect 175 2275 209 2751
rect -209 1557 -175 2033
rect -113 1557 -79 2033
rect -17 1557 17 2033
rect 79 1557 113 2033
rect 175 1557 209 2033
rect -209 839 -175 1315
rect -113 839 -79 1315
rect -17 839 17 1315
rect 79 839 113 1315
rect 175 839 209 1315
rect -209 121 -175 597
rect -113 121 -79 597
rect -17 121 17 597
rect 79 121 113 597
rect 175 121 209 597
rect -209 -597 -175 -121
rect -113 -597 -79 -121
rect -17 -597 17 -121
rect 79 -597 113 -121
rect 175 -597 209 -121
rect -209 -1315 -175 -839
rect -113 -1315 -79 -839
rect -17 -1315 17 -839
rect 79 -1315 113 -839
rect 175 -1315 209 -839
rect -209 -2033 -175 -1557
rect -113 -2033 -79 -1557
rect -17 -2033 17 -1557
rect 79 -2033 113 -1557
rect 175 -2033 209 -1557
rect -209 -2751 -175 -2275
rect -113 -2751 -79 -2275
rect -17 -2751 17 -2275
rect 79 -2751 113 -2275
rect 175 -2751 209 -2275
<< psubdiff >>
rect -323 2903 -227 2937
rect 227 2903 323 2937
rect -323 2841 -289 2903
rect 289 2841 323 2903
rect -323 -2903 -289 -2841
rect 289 -2903 323 -2841
rect -323 -2937 -227 -2903
rect 227 -2937 323 -2903
<< psubdiffcont >>
rect -227 2903 227 2937
rect -323 -2841 -289 2841
rect 289 -2841 323 2841
rect -227 -2937 227 -2903
<< poly >>
rect -177 2835 -111 2851
rect -177 2801 -161 2835
rect -127 2801 -111 2835
rect -177 2785 -111 2801
rect 15 2835 81 2851
rect 15 2801 31 2835
rect 65 2801 81 2835
rect -159 2763 -129 2785
rect -63 2763 -33 2789
rect 15 2785 81 2801
rect 33 2763 63 2785
rect 129 2763 159 2789
rect -159 2237 -129 2263
rect -63 2241 -33 2263
rect -81 2225 -15 2241
rect 33 2237 63 2263
rect 129 2241 159 2263
rect -81 2191 -65 2225
rect -31 2191 -15 2225
rect -81 2175 -15 2191
rect 111 2225 177 2241
rect 111 2191 127 2225
rect 161 2191 177 2225
rect 111 2175 177 2191
rect -81 2117 -15 2133
rect -81 2083 -65 2117
rect -31 2083 -15 2117
rect -159 2045 -129 2071
rect -81 2067 -15 2083
rect 111 2117 177 2133
rect 111 2083 127 2117
rect 161 2083 177 2117
rect -63 2045 -33 2067
rect 33 2045 63 2071
rect 111 2067 177 2083
rect 129 2045 159 2067
rect -159 1523 -129 1545
rect -177 1507 -111 1523
rect -63 1519 -33 1545
rect 33 1523 63 1545
rect -177 1473 -161 1507
rect -127 1473 -111 1507
rect -177 1457 -111 1473
rect 15 1507 81 1523
rect 129 1519 159 1545
rect 15 1473 31 1507
rect 65 1473 81 1507
rect 15 1457 81 1473
rect -177 1399 -111 1415
rect -177 1365 -161 1399
rect -127 1365 -111 1399
rect -177 1349 -111 1365
rect 15 1399 81 1415
rect 15 1365 31 1399
rect 65 1365 81 1399
rect -159 1327 -129 1349
rect -63 1327 -33 1353
rect 15 1349 81 1365
rect 33 1327 63 1349
rect 129 1327 159 1353
rect -159 801 -129 827
rect -63 805 -33 827
rect -81 789 -15 805
rect 33 801 63 827
rect 129 805 159 827
rect -81 755 -65 789
rect -31 755 -15 789
rect -81 739 -15 755
rect 111 789 177 805
rect 111 755 127 789
rect 161 755 177 789
rect 111 739 177 755
rect -81 681 -15 697
rect -81 647 -65 681
rect -31 647 -15 681
rect -159 609 -129 635
rect -81 631 -15 647
rect 111 681 177 697
rect 111 647 127 681
rect 161 647 177 681
rect -63 609 -33 631
rect 33 609 63 635
rect 111 631 177 647
rect 129 609 159 631
rect -159 87 -129 109
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 33 -109 63 -87
rect 129 -109 159 -83
rect -159 -635 -129 -609
rect -63 -631 -33 -609
rect -81 -647 -15 -631
rect 33 -635 63 -609
rect 129 -631 159 -609
rect -81 -681 -65 -647
rect -31 -681 -15 -647
rect -81 -697 -15 -681
rect 111 -647 177 -631
rect 111 -681 127 -647
rect 161 -681 177 -647
rect 111 -697 177 -681
rect -81 -755 -15 -739
rect -81 -789 -65 -755
rect -31 -789 -15 -755
rect -159 -827 -129 -801
rect -81 -805 -15 -789
rect 111 -755 177 -739
rect 111 -789 127 -755
rect 161 -789 177 -755
rect -63 -827 -33 -805
rect 33 -827 63 -801
rect 111 -805 177 -789
rect 129 -827 159 -805
rect -159 -1349 -129 -1327
rect -177 -1365 -111 -1349
rect -63 -1353 -33 -1327
rect 33 -1349 63 -1327
rect -177 -1399 -161 -1365
rect -127 -1399 -111 -1365
rect -177 -1415 -111 -1399
rect 15 -1365 81 -1349
rect 129 -1353 159 -1327
rect 15 -1399 31 -1365
rect 65 -1399 81 -1365
rect 15 -1415 81 -1399
rect -177 -1473 -111 -1457
rect -177 -1507 -161 -1473
rect -127 -1507 -111 -1473
rect -177 -1523 -111 -1507
rect 15 -1473 81 -1457
rect 15 -1507 31 -1473
rect 65 -1507 81 -1473
rect -159 -1545 -129 -1523
rect -63 -1545 -33 -1519
rect 15 -1523 81 -1507
rect 33 -1545 63 -1523
rect 129 -1545 159 -1519
rect -159 -2071 -129 -2045
rect -63 -2067 -33 -2045
rect -81 -2083 -15 -2067
rect 33 -2071 63 -2045
rect 129 -2067 159 -2045
rect -81 -2117 -65 -2083
rect -31 -2117 -15 -2083
rect -81 -2133 -15 -2117
rect 111 -2083 177 -2067
rect 111 -2117 127 -2083
rect 161 -2117 177 -2083
rect 111 -2133 177 -2117
rect -81 -2191 -15 -2175
rect -81 -2225 -65 -2191
rect -31 -2225 -15 -2191
rect -159 -2263 -129 -2237
rect -81 -2241 -15 -2225
rect 111 -2191 177 -2175
rect 111 -2225 127 -2191
rect 161 -2225 177 -2191
rect -63 -2263 -33 -2241
rect 33 -2263 63 -2237
rect 111 -2241 177 -2225
rect 129 -2263 159 -2241
rect -159 -2785 -129 -2763
rect -177 -2801 -111 -2785
rect -63 -2789 -33 -2763
rect 33 -2785 63 -2763
rect -177 -2835 -161 -2801
rect -127 -2835 -111 -2801
rect -177 -2851 -111 -2835
rect 15 -2801 81 -2785
rect 129 -2789 159 -2763
rect 15 -2835 31 -2801
rect 65 -2835 81 -2801
rect 15 -2851 81 -2835
<< polycont >>
rect -161 2801 -127 2835
rect 31 2801 65 2835
rect -65 2191 -31 2225
rect 127 2191 161 2225
rect -65 2083 -31 2117
rect 127 2083 161 2117
rect -161 1473 -127 1507
rect 31 1473 65 1507
rect -161 1365 -127 1399
rect 31 1365 65 1399
rect -65 755 -31 789
rect 127 755 161 789
rect -65 647 -31 681
rect 127 647 161 681
rect -161 37 -127 71
rect 31 37 65 71
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect -65 -681 -31 -647
rect 127 -681 161 -647
rect -65 -789 -31 -755
rect 127 -789 161 -755
rect -161 -1399 -127 -1365
rect 31 -1399 65 -1365
rect -161 -1507 -127 -1473
rect 31 -1507 65 -1473
rect -65 -2117 -31 -2083
rect 127 -2117 161 -2083
rect -65 -2225 -31 -2191
rect 127 -2225 161 -2191
rect -161 -2835 -127 -2801
rect 31 -2835 65 -2801
<< locali >>
rect -323 2903 -227 2937
rect 227 2903 323 2937
rect -323 2841 -289 2903
rect 289 2841 323 2903
rect -177 2801 -161 2835
rect -127 2801 -111 2835
rect 15 2801 31 2835
rect 65 2801 81 2835
rect -209 2751 -175 2767
rect -209 2259 -175 2275
rect -113 2751 -79 2767
rect -113 2259 -79 2275
rect -17 2751 17 2767
rect -17 2259 17 2275
rect 79 2751 113 2767
rect 79 2259 113 2275
rect 175 2751 209 2767
rect 175 2259 209 2275
rect -81 2191 -65 2225
rect -31 2191 -15 2225
rect 111 2191 127 2225
rect 161 2191 177 2225
rect -81 2083 -65 2117
rect -31 2083 -15 2117
rect 111 2083 127 2117
rect 161 2083 177 2117
rect -209 2033 -175 2049
rect -209 1541 -175 1557
rect -113 2033 -79 2049
rect -113 1541 -79 1557
rect -17 2033 17 2049
rect -17 1541 17 1557
rect 79 2033 113 2049
rect 79 1541 113 1557
rect 175 2033 209 2049
rect 175 1541 209 1557
rect -177 1473 -161 1507
rect -127 1473 -111 1507
rect 15 1473 31 1507
rect 65 1473 81 1507
rect -177 1365 -161 1399
rect -127 1365 -111 1399
rect 15 1365 31 1399
rect 65 1365 81 1399
rect -209 1315 -175 1331
rect -209 823 -175 839
rect -113 1315 -79 1331
rect -113 823 -79 839
rect -17 1315 17 1331
rect -17 823 17 839
rect 79 1315 113 1331
rect 79 823 113 839
rect 175 1315 209 1331
rect 175 823 209 839
rect -81 755 -65 789
rect -31 755 -15 789
rect 111 755 127 789
rect 161 755 177 789
rect -81 647 -65 681
rect -31 647 -15 681
rect 111 647 127 681
rect 161 647 177 681
rect -209 597 -175 613
rect -209 105 -175 121
rect -113 597 -79 613
rect -113 105 -79 121
rect -17 597 17 613
rect -17 105 17 121
rect 79 597 113 613
rect 79 105 113 121
rect 175 597 209 613
rect 175 105 209 121
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -209 -121 -175 -105
rect -209 -613 -175 -597
rect -113 -121 -79 -105
rect -113 -613 -79 -597
rect -17 -121 17 -105
rect -17 -613 17 -597
rect 79 -121 113 -105
rect 79 -613 113 -597
rect 175 -121 209 -105
rect 175 -613 209 -597
rect -81 -681 -65 -647
rect -31 -681 -15 -647
rect 111 -681 127 -647
rect 161 -681 177 -647
rect -81 -789 -65 -755
rect -31 -789 -15 -755
rect 111 -789 127 -755
rect 161 -789 177 -755
rect -209 -839 -175 -823
rect -209 -1331 -175 -1315
rect -113 -839 -79 -823
rect -113 -1331 -79 -1315
rect -17 -839 17 -823
rect -17 -1331 17 -1315
rect 79 -839 113 -823
rect 79 -1331 113 -1315
rect 175 -839 209 -823
rect 175 -1331 209 -1315
rect -177 -1399 -161 -1365
rect -127 -1399 -111 -1365
rect 15 -1399 31 -1365
rect 65 -1399 81 -1365
rect -177 -1507 -161 -1473
rect -127 -1507 -111 -1473
rect 15 -1507 31 -1473
rect 65 -1507 81 -1473
rect -209 -1557 -175 -1541
rect -209 -2049 -175 -2033
rect -113 -1557 -79 -1541
rect -113 -2049 -79 -2033
rect -17 -1557 17 -1541
rect -17 -2049 17 -2033
rect 79 -1557 113 -1541
rect 79 -2049 113 -2033
rect 175 -1557 209 -1541
rect 175 -2049 209 -2033
rect -81 -2117 -65 -2083
rect -31 -2117 -15 -2083
rect 111 -2117 127 -2083
rect 161 -2117 177 -2083
rect -81 -2225 -65 -2191
rect -31 -2225 -15 -2191
rect 111 -2225 127 -2191
rect 161 -2225 177 -2191
rect -209 -2275 -175 -2259
rect -209 -2767 -175 -2751
rect -113 -2275 -79 -2259
rect -113 -2767 -79 -2751
rect -17 -2275 17 -2259
rect -17 -2767 17 -2751
rect 79 -2275 113 -2259
rect 79 -2767 113 -2751
rect 175 -2275 209 -2259
rect 175 -2767 209 -2751
rect -177 -2835 -161 -2801
rect -127 -2835 -111 -2801
rect 15 -2835 31 -2801
rect 65 -2835 81 -2801
rect -323 -2903 -289 -2841
rect 289 -2903 323 -2841
rect -323 -2937 -227 -2903
rect 227 -2937 323 -2903
<< viali >>
rect -161 2801 -127 2835
rect 31 2801 65 2835
rect -209 2275 -175 2751
rect -113 2275 -79 2751
rect -17 2275 17 2751
rect 79 2275 113 2751
rect 175 2275 209 2751
rect -65 2191 -31 2225
rect 127 2191 161 2225
rect -65 2083 -31 2117
rect 127 2083 161 2117
rect -209 1557 -175 2033
rect -113 1557 -79 2033
rect -17 1557 17 2033
rect 79 1557 113 2033
rect 175 1557 209 2033
rect -161 1473 -127 1507
rect 31 1473 65 1507
rect -161 1365 -127 1399
rect 31 1365 65 1399
rect -209 839 -175 1315
rect -113 839 -79 1315
rect -17 839 17 1315
rect 79 839 113 1315
rect 175 839 209 1315
rect -65 755 -31 789
rect 127 755 161 789
rect -65 647 -31 681
rect 127 647 161 681
rect -209 121 -175 597
rect -113 121 -79 597
rect -17 121 17 597
rect 79 121 113 597
rect 175 121 209 597
rect -161 37 -127 71
rect 31 37 65 71
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect -209 -597 -175 -121
rect -113 -597 -79 -121
rect -17 -597 17 -121
rect 79 -597 113 -121
rect 175 -597 209 -121
rect -65 -681 -31 -647
rect 127 -681 161 -647
rect -65 -789 -31 -755
rect 127 -789 161 -755
rect -209 -1315 -175 -839
rect -113 -1315 -79 -839
rect -17 -1315 17 -839
rect 79 -1315 113 -839
rect 175 -1315 209 -839
rect -161 -1399 -127 -1365
rect 31 -1399 65 -1365
rect -161 -1507 -127 -1473
rect 31 -1507 65 -1473
rect -209 -2033 -175 -1557
rect -113 -2033 -79 -1557
rect -17 -2033 17 -1557
rect 79 -2033 113 -1557
rect 175 -2033 209 -1557
rect -65 -2117 -31 -2083
rect 127 -2117 161 -2083
rect -65 -2225 -31 -2191
rect 127 -2225 161 -2191
rect -209 -2751 -175 -2275
rect -113 -2751 -79 -2275
rect -17 -2751 17 -2275
rect 79 -2751 113 -2275
rect 175 -2751 209 -2275
rect -161 -2835 -127 -2801
rect 31 -2835 65 -2801
<< metal1 >>
rect -173 2835 -115 2841
rect -173 2801 -161 2835
rect -127 2801 -115 2835
rect -173 2795 -115 2801
rect 19 2835 77 2841
rect 19 2801 31 2835
rect 65 2801 77 2835
rect 19 2795 77 2801
rect -215 2751 -169 2763
rect -215 2275 -209 2751
rect -175 2275 -169 2751
rect -215 2263 -169 2275
rect -119 2751 -73 2763
rect -119 2275 -113 2751
rect -79 2275 -73 2751
rect -119 2263 -73 2275
rect -23 2751 23 2763
rect -23 2275 -17 2751
rect 17 2275 23 2751
rect -23 2263 23 2275
rect 73 2751 119 2763
rect 73 2275 79 2751
rect 113 2275 119 2751
rect 73 2263 119 2275
rect 169 2751 215 2763
rect 169 2275 175 2751
rect 209 2275 215 2751
rect 169 2263 215 2275
rect -77 2225 -19 2231
rect -77 2191 -65 2225
rect -31 2191 -19 2225
rect -77 2185 -19 2191
rect 115 2225 173 2231
rect 115 2191 127 2225
rect 161 2191 173 2225
rect 115 2185 173 2191
rect -77 2117 -19 2123
rect -77 2083 -65 2117
rect -31 2083 -19 2117
rect -77 2077 -19 2083
rect 115 2117 173 2123
rect 115 2083 127 2117
rect 161 2083 173 2117
rect 115 2077 173 2083
rect -215 2033 -169 2045
rect -215 1557 -209 2033
rect -175 1557 -169 2033
rect -215 1545 -169 1557
rect -119 2033 -73 2045
rect -119 1557 -113 2033
rect -79 1557 -73 2033
rect -119 1545 -73 1557
rect -23 2033 23 2045
rect -23 1557 -17 2033
rect 17 1557 23 2033
rect -23 1545 23 1557
rect 73 2033 119 2045
rect 73 1557 79 2033
rect 113 1557 119 2033
rect 73 1545 119 1557
rect 169 2033 215 2045
rect 169 1557 175 2033
rect 209 1557 215 2033
rect 169 1545 215 1557
rect -173 1507 -115 1513
rect -173 1473 -161 1507
rect -127 1473 -115 1507
rect -173 1467 -115 1473
rect 19 1507 77 1513
rect 19 1473 31 1507
rect 65 1473 77 1507
rect 19 1467 77 1473
rect -173 1399 -115 1405
rect -173 1365 -161 1399
rect -127 1365 -115 1399
rect -173 1359 -115 1365
rect 19 1399 77 1405
rect 19 1365 31 1399
rect 65 1365 77 1399
rect 19 1359 77 1365
rect -215 1315 -169 1327
rect -215 839 -209 1315
rect -175 839 -169 1315
rect -215 827 -169 839
rect -119 1315 -73 1327
rect -119 839 -113 1315
rect -79 839 -73 1315
rect -119 827 -73 839
rect -23 1315 23 1327
rect -23 839 -17 1315
rect 17 839 23 1315
rect -23 827 23 839
rect 73 1315 119 1327
rect 73 839 79 1315
rect 113 839 119 1315
rect 73 827 119 839
rect 169 1315 215 1327
rect 169 839 175 1315
rect 209 839 215 1315
rect 169 827 215 839
rect -77 789 -19 795
rect -77 755 -65 789
rect -31 755 -19 789
rect -77 749 -19 755
rect 115 789 173 795
rect 115 755 127 789
rect 161 755 173 789
rect 115 749 173 755
rect -77 681 -19 687
rect -77 647 -65 681
rect -31 647 -19 681
rect -77 641 -19 647
rect 115 681 173 687
rect 115 647 127 681
rect 161 647 173 681
rect 115 641 173 647
rect -215 597 -169 609
rect -215 121 -209 597
rect -175 121 -169 597
rect -215 109 -169 121
rect -119 597 -73 609
rect -119 121 -113 597
rect -79 121 -73 597
rect -119 109 -73 121
rect -23 597 23 609
rect -23 121 -17 597
rect 17 121 23 597
rect -23 109 23 121
rect 73 597 119 609
rect 73 121 79 597
rect 113 121 119 597
rect 73 109 119 121
rect 169 597 215 609
rect 169 121 175 597
rect 209 121 215 597
rect 169 109 215 121
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect -215 -121 -169 -109
rect -215 -597 -209 -121
rect -175 -597 -169 -121
rect -215 -609 -169 -597
rect -119 -121 -73 -109
rect -119 -597 -113 -121
rect -79 -597 -73 -121
rect -119 -609 -73 -597
rect -23 -121 23 -109
rect -23 -597 -17 -121
rect 17 -597 23 -121
rect -23 -609 23 -597
rect 73 -121 119 -109
rect 73 -597 79 -121
rect 113 -597 119 -121
rect 73 -609 119 -597
rect 169 -121 215 -109
rect 169 -597 175 -121
rect 209 -597 215 -121
rect 169 -609 215 -597
rect -77 -647 -19 -641
rect -77 -681 -65 -647
rect -31 -681 -19 -647
rect -77 -687 -19 -681
rect 115 -647 173 -641
rect 115 -681 127 -647
rect 161 -681 173 -647
rect 115 -687 173 -681
rect -77 -755 -19 -749
rect -77 -789 -65 -755
rect -31 -789 -19 -755
rect -77 -795 -19 -789
rect 115 -755 173 -749
rect 115 -789 127 -755
rect 161 -789 173 -755
rect 115 -795 173 -789
rect -215 -839 -169 -827
rect -215 -1315 -209 -839
rect -175 -1315 -169 -839
rect -215 -1327 -169 -1315
rect -119 -839 -73 -827
rect -119 -1315 -113 -839
rect -79 -1315 -73 -839
rect -119 -1327 -73 -1315
rect -23 -839 23 -827
rect -23 -1315 -17 -839
rect 17 -1315 23 -839
rect -23 -1327 23 -1315
rect 73 -839 119 -827
rect 73 -1315 79 -839
rect 113 -1315 119 -839
rect 73 -1327 119 -1315
rect 169 -839 215 -827
rect 169 -1315 175 -839
rect 209 -1315 215 -839
rect 169 -1327 215 -1315
rect -173 -1365 -115 -1359
rect -173 -1399 -161 -1365
rect -127 -1399 -115 -1365
rect -173 -1405 -115 -1399
rect 19 -1365 77 -1359
rect 19 -1399 31 -1365
rect 65 -1399 77 -1365
rect 19 -1405 77 -1399
rect -173 -1473 -115 -1467
rect -173 -1507 -161 -1473
rect -127 -1507 -115 -1473
rect -173 -1513 -115 -1507
rect 19 -1473 77 -1467
rect 19 -1507 31 -1473
rect 65 -1507 77 -1473
rect 19 -1513 77 -1507
rect -215 -1557 -169 -1545
rect -215 -2033 -209 -1557
rect -175 -2033 -169 -1557
rect -215 -2045 -169 -2033
rect -119 -1557 -73 -1545
rect -119 -2033 -113 -1557
rect -79 -2033 -73 -1557
rect -119 -2045 -73 -2033
rect -23 -1557 23 -1545
rect -23 -2033 -17 -1557
rect 17 -2033 23 -1557
rect -23 -2045 23 -2033
rect 73 -1557 119 -1545
rect 73 -2033 79 -1557
rect 113 -2033 119 -1557
rect 73 -2045 119 -2033
rect 169 -1557 215 -1545
rect 169 -2033 175 -1557
rect 209 -2033 215 -1557
rect 169 -2045 215 -2033
rect -77 -2083 -19 -2077
rect -77 -2117 -65 -2083
rect -31 -2117 -19 -2083
rect -77 -2123 -19 -2117
rect 115 -2083 173 -2077
rect 115 -2117 127 -2083
rect 161 -2117 173 -2083
rect 115 -2123 173 -2117
rect -77 -2191 -19 -2185
rect -77 -2225 -65 -2191
rect -31 -2225 -19 -2191
rect -77 -2231 -19 -2225
rect 115 -2191 173 -2185
rect 115 -2225 127 -2191
rect 161 -2225 173 -2191
rect 115 -2231 173 -2225
rect -215 -2275 -169 -2263
rect -215 -2751 -209 -2275
rect -175 -2751 -169 -2275
rect -215 -2763 -169 -2751
rect -119 -2275 -73 -2263
rect -119 -2751 -113 -2275
rect -79 -2751 -73 -2275
rect -119 -2763 -73 -2751
rect -23 -2275 23 -2263
rect -23 -2751 -17 -2275
rect 17 -2751 23 -2275
rect -23 -2763 23 -2751
rect 73 -2275 119 -2263
rect 73 -2751 79 -2275
rect 113 -2751 119 -2275
rect 73 -2763 119 -2751
rect 169 -2275 215 -2263
rect 169 -2751 175 -2275
rect 209 -2751 215 -2275
rect 169 -2763 215 -2751
rect -173 -2801 -115 -2795
rect -173 -2835 -161 -2801
rect -127 -2835 -115 -2801
rect -173 -2841 -115 -2835
rect 19 -2801 77 -2795
rect 19 -2835 31 -2801
rect 65 -2835 77 -2801
rect 19 -2841 77 -2835
<< properties >>
string FIXED_BBOX -306 -2920 306 2920
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 8 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
