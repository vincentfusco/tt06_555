magic
tech sky130A
magscale 1 2
timestamp 1711057506
<< error_p >>
rect 26831 28007 26866 28041
rect 26832 27988 26866 28007
rect 26640 27939 26702 27945
rect 26640 27905 26652 27939
rect 26640 27899 26702 27905
rect 26640 25811 26702 25817
rect 26640 25777 26652 25811
rect 26640 25771 26702 25777
rect 26640 25703 26702 25709
rect 26640 25669 26652 25703
rect 26640 25663 26702 25669
rect 26640 23575 26702 23581
rect 26640 23541 26652 23575
rect 26640 23535 26702 23541
rect 26640 23467 26702 23473
rect 26640 23433 26652 23467
rect 26640 23427 26702 23433
rect 26640 21339 26702 21345
rect 26640 21305 26652 21339
rect 26640 21299 26702 21305
rect 26640 21231 26702 21237
rect 26640 21197 26652 21231
rect 26640 21191 26702 21197
rect 11400 19292 11446 19304
rect 11928 19292 11974 19304
rect 11400 19258 11406 19292
rect 11928 19258 11934 19292
rect 11400 19246 11446 19258
rect 11928 19246 11974 19258
rect 26640 19103 26702 19109
rect 26640 19069 26652 19103
rect 26640 19063 26702 19069
rect 11400 18976 11446 18988
rect 11928 18976 11974 18988
rect 11400 18942 11406 18976
rect 11928 18942 11934 18976
rect 26851 18967 26866 27988
rect 26885 27954 26920 27988
rect 26885 18967 26919 27954
rect 27049 27886 27111 27892
rect 27049 27852 27061 27886
rect 27049 27846 27111 27852
rect 27049 25758 27111 25764
rect 27049 25724 27061 25758
rect 27049 25718 27111 25724
rect 27049 25650 27111 25656
rect 27049 25616 27061 25650
rect 27049 25610 27111 25616
rect 27049 23522 27111 23528
rect 27049 23488 27061 23522
rect 27049 23482 27111 23488
rect 27049 23414 27111 23420
rect 27049 23380 27061 23414
rect 27049 23374 27111 23380
rect 27049 21286 27111 21292
rect 27049 21252 27061 21286
rect 27049 21246 27111 21252
rect 27049 21178 27111 21184
rect 27049 21144 27061 21178
rect 27049 21138 27111 21144
rect 27867 20178 28319 20210
rect 27867 20144 28319 20156
rect 29450 20118 29484 20136
rect 27241 20045 27275 20063
rect 27241 20009 27311 20045
rect 27258 19975 27329 20009
rect 27049 19050 27111 19056
rect 27049 19016 27061 19050
rect 27049 19010 27111 19016
rect 11400 18930 11446 18942
rect 11928 18930 11974 18942
rect 26885 18933 26900 18967
rect 27258 18914 27328 19975
rect 27258 18878 27311 18914
rect 27799 18861 27814 20009
rect 27833 18861 27867 20060
rect 28945 20048 29397 20080
rect 28945 20014 29397 20026
rect 28319 19879 28353 19933
rect 27833 18827 27848 18861
rect 28338 18784 28353 19879
rect 28372 19845 28407 19879
rect 28372 18784 28406 19845
rect 28372 18750 28387 18784
rect 28877 18731 28892 19879
rect 28911 18731 28945 19930
rect 28911 18697 28926 18731
rect 29414 18654 29484 20118
rect 29936 19988 29970 20006
rect 29936 19952 30006 19988
rect 29953 19950 30024 19952
rect 29953 19929 30475 19950
rect 29953 19918 30509 19929
rect 29953 19896 30023 19918
rect 30475 19896 30509 19918
rect 31067 19911 31101 19929
rect 29953 19884 30509 19896
rect 29953 19862 30024 19884
rect 30474 19875 30509 19884
rect 29414 18618 29467 18654
rect 29953 18601 30023 19862
rect 29953 18565 30006 18601
rect 11500 18518 11546 18530
rect 11810 18518 11856 18530
rect 30494 18524 30509 19875
rect 30528 19873 30563 19875
rect 30528 19841 31014 19873
rect 30528 19819 30562 19841
rect 30528 19807 31014 19819
rect 30528 19785 30563 19807
rect 30528 18524 30562 19785
rect 11500 18484 11506 18518
rect 11810 18484 11816 18518
rect 30528 18490 30543 18524
rect 11500 18472 11546 18484
rect 11810 18472 11856 18484
rect 31031 18447 31101 19911
rect 31031 18411 31084 18447
rect 11500 18202 11546 18214
rect 11810 18202 11856 18214
rect 11500 18168 11506 18202
rect 11810 18168 11816 18202
rect 11500 18156 11546 18168
rect 11810 18156 11856 18168
rect 4726 14974 4772 14986
rect 5254 14974 5300 14986
rect 4726 14940 4732 14974
rect 5254 14940 5260 14974
rect 4726 14928 4772 14940
rect 5254 14928 5300 14940
rect 4726 14658 4772 14670
rect 5254 14658 5300 14670
rect 4726 14624 4732 14658
rect 5254 14624 5260 14658
rect 4726 14612 4772 14624
rect 5254 14612 5300 14624
rect 4826 14200 4872 14212
rect 5136 14200 5182 14212
rect 4826 14166 4832 14200
rect 5136 14166 5142 14200
rect 4826 14154 4872 14166
rect 5136 14154 5182 14166
rect 4826 13884 4872 13896
rect 5136 13884 5182 13896
rect 4826 13850 4832 13884
rect 5136 13850 5142 13884
rect 4826 13838 4872 13850
rect 5136 13838 5182 13850
rect 24246 4892 24308 4898
rect 24246 4858 24258 4892
rect 24246 4852 24308 4858
rect 24246 3782 24308 3788
rect 24246 3748 24258 3782
rect 24246 3742 24308 3748
rect 24246 3674 24308 3680
rect 24246 3640 24258 3674
rect 24246 3634 24308 3640
rect 24246 2564 24308 2570
rect 24246 2530 24258 2564
rect 24246 2524 24308 2530
rect 24246 2456 24308 2462
rect 24246 2422 24258 2456
rect 24246 2416 24308 2422
rect 24246 1346 24308 1352
rect 24246 1312 24258 1346
rect 24246 1306 24308 1312
rect 24246 1238 24308 1244
rect 24246 1204 24258 1238
rect 24246 1198 24308 1204
rect 24246 128 24308 134
rect 24246 94 24258 128
rect 24246 88 24308 94
<< error_s >>
rect 8493 3459 8714 3469
rect 8747 2831 8968 3459
rect 9148 2421 9169 3227
rect 9176 2821 9423 3459
rect 9176 2393 9197 2821
rect 9577 2421 9598 3227
rect 9605 2821 9852 3459
rect 9605 2393 9626 2821
rect 10006 2421 10027 3227
rect 10034 2821 10281 3459
rect 10034 2393 10055 2821
rect 10435 2421 10456 3227
rect 10463 2821 10710 3459
rect 10463 2393 10484 2821
rect 10864 2421 10885 3227
rect 10892 2821 11139 3459
rect 10892 2393 10913 2821
rect 17565 1811 17599 1829
rect 17529 352 17599 1811
rect 17529 347 17600 352
rect 17529 311 17582 347
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use comp_n  X_COMP_N
timestamp 1711057506
transform 1 0 29431 0 1 4920
box 18500 1578 24043 5238
use comp_p  X_COMP_P1
timestamp 1711053111
transform 1 0 26493 0 1 18384
box -53 -2000 5669 9693
use inv  X_INV1
timestamp 1711045747
transform 1 0 8352 0 1 1649
box -60 547 369 1820
use inv  X_INV2[0]
timestamp 1711045747
transform 1 0 9236 0 1 1639
box -60 547 369 1820
use inv  X_INV2[1]
timestamp 1711045747
transform 1 0 8807 0 1 1639
box -60 547 369 1820
use inv  X_INV3[0]
timestamp 1711045747
transform 1 0 10952 0 1 1639
box -60 547 369 1820
use inv  X_INV3[1]
timestamp 1711045747
transform 1 0 10523 0 1 1639
box -60 547 369 1820
use inv  X_INV3[2]
timestamp 1711045747
transform 1 0 10094 0 1 1639
box -60 547 369 1820
use inv  X_INV3[3]
timestamp 1711045747
transform 1 0 9665 0 1 1639
box -60 547 369 1820
use sr_latch  X_SR_LATCH
timestamp 1711045747
transform 1 0 8745 0 1 14056
box -4457 -2000 3703 5706
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_bias
timestamp 1711041810
transform 1 0 17286 0 1 1045
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_44Y62X  XMn_discharge
timestamp 1711041017
transform 1 0 24277 0 1 2493
box -231 -2537 2431 2537
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_bias
timestamp 1711036998
transform 1 0 17825 0 1 1501
box -296 -1219 296 1219
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_1
timestamp 1711037431
transform 1 0 10561 0 1 -2770
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_2
timestamp 1711037431
transform 1 0 13413 0 1 -2446
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_3
timestamp 1711037431
transform 1 0 14119 0 1 -2418
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_4
timestamp 1711037431
transform 1 0 14973 0 1 -2418
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bot
timestamp 1711037431
transform 1 0 9795 0 1 -2828
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_mid
timestamp 1711037431
transform 1 0 9089 0 1 -2946
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_top
timestamp 1711037431
transform 1 0 8383 0 1 -2976
box -307 -1282 307 1282
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 DO_OUT
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 V_DISCH_O
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 V_THRESH_I
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 V_TRIG_B_I
port 5 nsew
<< end >>
