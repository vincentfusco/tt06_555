** sch_path: /home/vincef/projects/tt06_555/xsch/ip/comparators/comp_p.sch
.subckt comp_p vinp vout vdd vss vinn vbias_p
*.PININFO vdd:B vss:B vbias_p:I vinn:I vinp:I vout:O
XMp_inn1 latch_left vinn tail vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 m=4
XMp_inp1 latch_right vinp tail vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 m=4
XMn_diode_left1 latch_left latch_left vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XMn_cs_left latch_right latch_left vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=1
XMn_diode_right latch_right latch_right vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XMn_cs_right1 latch_left latch_right vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=1
XMp_tail tail vbias_p vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=10 nf=1 m=1
XMn_out_right vout latch_right vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=1
XMn_out_left out_left latch_left vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=1
XMp_diode_left1 out_left out_left vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 m=1
XMp_out vout out_left vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 m=1
.ends
.end
