magic
tech sky130A
timestamp 1712095588
<< metal2 >>
rect 2352 5628 3724 6076
rect 2660 5600 3416 5628
rect 1652 5572 1876 5600
rect 1596 5544 1904 5572
rect 1540 5516 1932 5544
rect 1484 5488 1960 5516
rect 1456 5460 1988 5488
rect 1400 5432 1988 5460
rect 1372 5404 2016 5432
rect 1316 5376 2044 5404
rect 1288 5348 2044 5376
rect 1288 5320 2072 5348
rect 1260 5292 2072 5320
rect 1260 5236 2100 5292
rect 2688 5236 3388 5600
rect 4228 5572 4452 5600
rect 4172 5544 4480 5572
rect 4144 5516 4536 5544
rect 4116 5488 4592 5516
rect 4116 5460 4620 5488
rect 4088 5432 4676 5460
rect 4060 5404 4732 5432
rect 4060 5376 4760 5404
rect 4032 5348 4788 5376
rect 4004 5320 4788 5348
rect 4004 5292 4816 5320
rect 3976 5264 4816 5292
rect 3976 5236 4844 5264
rect 1260 5208 2044 5236
rect 2688 5208 3416 5236
rect 4032 5208 4844 5236
rect 1232 5180 2016 5208
rect 2604 5180 3500 5208
rect 4060 5180 4844 5208
rect 1260 5124 1988 5180
rect 2464 5152 3612 5180
rect 4116 5152 4844 5180
rect 2352 5124 3724 5152
rect 1260 5096 2016 5124
rect 2268 5096 3808 5124
rect 4088 5096 4816 5152
rect 1288 5068 2016 5096
rect 2184 5068 3892 5096
rect 4060 5068 4816 5096
rect 1288 5040 2044 5068
rect 2128 5040 3976 5068
rect 4032 5040 4788 5068
rect 1316 4984 4760 5040
rect 1344 4956 4732 4984
rect 1372 4928 4732 4956
rect 1372 4900 1540 4928
rect 1568 4900 4508 4928
rect 4536 4900 4704 4928
rect 1400 4872 1512 4900
rect 1400 4844 1456 4872
rect 1596 4844 4480 4900
rect 4592 4872 4676 4900
rect 4620 4844 4676 4872
rect 1624 4788 4452 4844
rect 1624 4760 2912 4788
rect 3164 4760 4480 4788
rect 1568 4732 2688 4760
rect 3388 4732 4508 4760
rect 1540 4704 2548 4732
rect 3528 4704 4536 4732
rect 1512 4676 2464 4704
rect 3640 4676 4592 4704
rect 1456 4648 2380 4676
rect 3724 4648 4620 4676
rect 1428 4620 2296 4648
rect 3780 4620 4648 4648
rect 1400 4592 2240 4620
rect 3864 4592 4676 4620
rect 1372 4564 2184 4592
rect 3920 4564 4704 4592
rect 1344 4536 2128 4564
rect 3976 4536 4732 4564
rect 1316 4508 2072 4536
rect 4004 4508 4760 4536
rect 1288 4480 2016 4508
rect 1260 4452 1960 4480
rect 1232 4424 1932 4452
rect 1204 4396 1876 4424
rect 1176 4368 1848 4396
rect 1148 4340 1820 4368
rect 1148 4312 1792 4340
rect 2240 4312 2324 4340
rect 1120 4284 1736 4312
rect 2184 4284 2352 4312
rect 1092 4256 1708 4284
rect 2156 4256 2352 4284
rect 1064 4228 1680 4256
rect 2156 4228 2380 4256
rect 1064 4200 1652 4228
rect 2184 4200 2380 4228
rect 1036 4172 1624 4200
rect 2184 4172 2408 4200
rect 1008 4144 1596 4172
rect 2212 4144 2408 4172
rect 1008 4116 1568 4144
rect 2212 4116 2436 4144
rect 980 4088 1540 4116
rect 2240 4088 2436 4116
rect 952 4032 1512 4088
rect 2240 4060 2464 4088
rect 2268 4032 2464 4060
rect 924 4004 1484 4032
rect 924 3976 1456 4004
rect 2296 3976 2492 4032
rect 896 3948 1428 3976
rect 868 3920 1428 3948
rect 2324 3948 2464 3976
rect 2324 3920 2408 3948
rect 868 3892 1400 3920
rect 2352 3892 2380 3920
rect 840 3836 1372 3892
rect 812 3808 1344 3836
rect 2940 3808 3136 4508
rect 4060 4480 4788 4508
rect 4116 4452 4816 4480
rect 4144 4424 4844 4452
rect 4200 4396 4872 4424
rect 4228 4368 4900 4396
rect 4256 4340 4928 4368
rect 3752 4312 3836 4340
rect 4312 4312 4956 4340
rect 3752 4284 3892 4312
rect 4340 4284 4956 4312
rect 3724 4228 3920 4284
rect 4368 4256 4984 4284
rect 4396 4228 5012 4256
rect 3696 4172 3892 4228
rect 4424 4200 5040 4228
rect 4452 4172 5040 4200
rect 3668 4144 3864 4172
rect 4480 4144 5068 4172
rect 3640 4116 3864 4144
rect 4508 4116 5096 4144
rect 3640 4088 3836 4116
rect 4536 4088 5096 4116
rect 3612 4060 3836 4088
rect 4564 4060 5124 4088
rect 3612 4032 3808 4060
rect 3584 4004 3808 4032
rect 4592 4004 5152 4060
rect 3584 3976 3780 4004
rect 4620 3976 5180 4004
rect 3612 3948 3780 3976
rect 4648 3948 5180 3976
rect 3668 3920 3752 3948
rect 4676 3892 5208 3948
rect 4704 3864 5236 3892
rect 4732 3836 5236 3864
rect 4732 3808 5264 3836
rect 812 3752 1316 3808
rect 2968 3780 3136 3808
rect 4760 3780 5264 3808
rect 1624 3752 1680 3780
rect 4396 3752 4480 3780
rect 4760 3752 5292 3780
rect 784 3696 1288 3752
rect 1596 3724 1736 3752
rect 4340 3724 4480 3752
rect 4788 3724 5292 3752
rect 1568 3696 1764 3724
rect 4312 3696 4508 3724
rect 756 3640 1260 3696
rect 1568 3668 1820 3696
rect 4256 3668 4508 3696
rect 4816 3668 5320 3724
rect 1540 3640 1848 3668
rect 4228 3640 4536 3668
rect 4844 3640 5320 3668
rect 756 3612 1232 3640
rect 1568 3612 1904 3640
rect 4172 3612 4508 3640
rect 728 3584 1232 3612
rect 1624 3584 1960 3612
rect 4144 3584 4480 3612
rect 4844 3584 5348 3640
rect 728 3528 1204 3584
rect 1652 3556 1988 3584
rect 4088 3556 4424 3584
rect 4872 3556 5348 3584
rect 1708 3528 1988 3556
rect 4116 3528 4396 3556
rect 4872 3528 5376 3556
rect 700 3500 1204 3528
rect 1736 3500 1960 3528
rect 4116 3500 4340 3528
rect 700 3444 1176 3500
rect 1792 3472 1932 3500
rect 1820 3444 1932 3472
rect 4144 3472 4284 3500
rect 4900 3472 5376 3528
rect 4144 3444 4256 3472
rect 4900 3444 5404 3472
rect 672 3360 1148 3444
rect 1876 3416 1904 3444
rect 4172 3416 4200 3444
rect 4928 3360 5404 3444
rect 672 3332 1120 3360
rect 644 3248 1120 3332
rect 4956 3276 5432 3360
rect 644 3192 1092 3248
rect 616 3108 1092 3192
rect 4984 3220 5432 3276
rect 2212 3108 2604 3164
rect 2828 3108 3220 3164
rect 3444 3108 3836 3164
rect 4984 3136 5460 3220
rect 616 2940 1064 3108
rect 2184 2996 2604 3108
rect 2800 2996 3220 3108
rect 3416 2996 3836 3108
rect 5012 3024 5460 3136
rect 2184 2940 2324 2996
rect 2800 2940 2940 2996
rect 3416 2940 3556 2996
rect 588 2632 1064 2940
rect 1316 2688 2044 2884
rect 2156 2856 2296 2940
rect 2324 2856 2492 2884
rect 2772 2856 2912 2940
rect 2940 2856 3108 2884
rect 3388 2856 3528 2940
rect 5012 2884 5488 3024
rect 3556 2856 3724 2884
rect 2156 2828 2548 2856
rect 2772 2828 3164 2856
rect 3388 2828 3780 2856
rect 2156 2800 2576 2828
rect 2772 2800 3192 2828
rect 3388 2800 3808 2828
rect 2156 2772 2604 2800
rect 2772 2772 3220 2800
rect 3388 2772 3836 2800
rect 2128 2744 2604 2772
rect 2744 2744 3220 2772
rect 3360 2744 3836 2772
rect 2128 2716 2296 2744
rect 2436 2716 2632 2744
rect 2744 2716 2912 2744
rect 3052 2716 3248 2744
rect 3360 2716 3528 2744
rect 3668 2716 3864 2744
rect 4032 2716 4760 2884
rect 5040 2716 5488 2884
rect 2156 2688 2268 2716
rect 2464 2688 2632 2716
rect 2772 2688 2884 2716
rect 3080 2688 3248 2716
rect 3388 2688 3500 2716
rect 3696 2688 3864 2716
rect 4060 2688 4760 2716
rect 616 2492 1064 2632
rect 2156 2576 2268 2604
rect 2128 2548 2268 2576
rect 2492 2548 2632 2688
rect 2772 2576 2884 2604
rect 2128 2520 2296 2548
rect 2464 2520 2632 2548
rect 2128 2492 2324 2520
rect 2436 2492 2632 2520
rect 2744 2548 2884 2576
rect 3108 2548 3248 2688
rect 3388 2576 3500 2604
rect 2744 2520 2912 2548
rect 3080 2520 3248 2548
rect 2744 2492 2940 2520
rect 3052 2492 3248 2520
rect 3360 2548 3500 2576
rect 3724 2548 3864 2688
rect 3360 2520 3528 2548
rect 3696 2520 3864 2548
rect 3360 2492 3556 2520
rect 3668 2492 3864 2520
rect 5012 2548 5488 2716
rect 616 2380 1092 2492
rect 2156 2464 2604 2492
rect 2772 2464 3220 2492
rect 3388 2464 3836 2492
rect 2156 2436 2576 2464
rect 2772 2436 3192 2464
rect 3388 2436 3808 2464
rect 5012 2436 5460 2548
rect 2184 2408 2548 2436
rect 2800 2408 3164 2436
rect 3416 2408 3780 2436
rect 2212 2380 2520 2408
rect 2828 2380 3136 2408
rect 3444 2380 3752 2408
rect 644 2352 1092 2380
rect 2268 2352 2464 2380
rect 2884 2352 3080 2380
rect 3500 2352 3696 2380
rect 4984 2352 5460 2436
rect 644 2240 1120 2352
rect 4984 2324 5432 2352
rect 672 2156 1148 2240
rect 4956 2212 5432 2324
rect 672 2128 1176 2156
rect 1848 2128 1904 2156
rect 4172 2128 4228 2156
rect 4928 2128 5404 2212
rect 700 2072 1176 2128
rect 1820 2100 1932 2128
rect 4144 2100 4256 2128
rect 4900 2100 5404 2128
rect 1764 2072 1960 2100
rect 4144 2072 4312 2100
rect 700 2044 1204 2072
rect 1736 2044 1960 2072
rect 4116 2044 4340 2072
rect 4900 2044 5376 2100
rect 728 1988 1204 2044
rect 1680 2016 1988 2044
rect 4088 2016 4396 2044
rect 4872 2016 5376 2044
rect 1652 1988 1988 2016
rect 4116 1988 4452 2016
rect 4872 1988 5348 2016
rect 728 1960 1232 1988
rect 1596 1960 1932 1988
rect 4144 1960 4480 1988
rect 756 1932 1232 1960
rect 1540 1932 1876 1960
rect 4200 1932 4536 1960
rect 4844 1932 5348 1988
rect 756 1876 1260 1932
rect 1540 1904 1848 1932
rect 4228 1904 4536 1932
rect 1568 1876 1792 1904
rect 4284 1876 4508 1904
rect 4816 1876 5320 1932
rect 784 1820 1288 1876
rect 1596 1848 1764 1876
rect 4312 1848 4508 1876
rect 1596 1820 1708 1848
rect 4368 1820 4480 1848
rect 4788 1820 5292 1876
rect 812 1792 1316 1820
rect 1624 1792 1680 1820
rect 4424 1792 4452 1820
rect 4760 1792 5292 1820
rect 812 1764 1344 1792
rect 840 1736 1344 1764
rect 840 1708 1372 1736
rect 868 1680 1372 1708
rect 868 1652 1400 1680
rect 2324 1652 2380 1680
rect 896 1624 1428 1652
rect 2324 1624 2436 1652
rect 896 1596 1456 1624
rect 924 1568 1456 1596
rect 2296 1568 2492 1624
rect 924 1540 1484 1568
rect 2268 1540 2492 1568
rect 952 1512 1512 1540
rect 2268 1512 2464 1540
rect 980 1484 1540 1512
rect 2240 1484 2464 1512
rect 980 1456 1568 1484
rect 2240 1456 2436 1484
rect 1008 1400 1596 1456
rect 2212 1428 2436 1456
rect 2212 1400 2408 1428
rect 1036 1372 1624 1400
rect 1064 1344 1652 1372
rect 2184 1344 2380 1400
rect 1092 1316 1708 1344
rect 1092 1288 1736 1316
rect 2156 1288 2352 1344
rect 1120 1260 1764 1288
rect 2212 1260 2324 1288
rect 1148 1232 1792 1260
rect 2268 1232 2324 1260
rect 1176 1204 1820 1232
rect 1204 1176 1876 1204
rect 1232 1148 1904 1176
rect 1232 1120 1932 1148
rect 1260 1092 1988 1120
rect 1288 1064 2044 1092
rect 2940 1064 3136 1792
rect 4760 1764 5264 1792
rect 4732 1736 5264 1764
rect 4704 1680 5236 1736
rect 3696 1652 3752 1680
rect 4676 1652 5208 1680
rect 3640 1624 3752 1652
rect 4648 1624 5208 1652
rect 3584 1568 3780 1624
rect 4648 1596 5180 1624
rect 4620 1568 5152 1596
rect 3612 1512 3808 1568
rect 4592 1540 5152 1568
rect 4564 1512 5124 1540
rect 3640 1456 3836 1512
rect 4536 1484 5124 1512
rect 4536 1456 5096 1484
rect 3668 1428 3864 1456
rect 4508 1428 5068 1456
rect 3668 1400 3892 1428
rect 4480 1400 5068 1428
rect 3696 1372 3892 1400
rect 4452 1372 5040 1400
rect 3696 1344 3920 1372
rect 4424 1344 5012 1372
rect 3724 1288 3920 1344
rect 4396 1316 5012 1344
rect 4368 1288 4984 1316
rect 3752 1260 3864 1288
rect 4312 1260 4956 1288
rect 3752 1232 3808 1260
rect 4284 1232 4928 1260
rect 4256 1204 4900 1232
rect 4228 1176 4900 1204
rect 4172 1148 4872 1176
rect 4144 1120 4844 1148
rect 4088 1092 4816 1120
rect 4060 1064 4788 1092
rect 1316 1036 2072 1064
rect 4004 1036 4760 1064
rect 1344 1008 2128 1036
rect 3948 1008 4732 1036
rect 1372 980 2184 1008
rect 3892 980 4704 1008
rect 1428 952 2240 980
rect 3836 952 4676 980
rect 1456 924 2324 952
rect 3752 924 4648 952
rect 1484 896 2408 924
rect 3696 896 4592 924
rect 1512 868 2492 896
rect 3584 868 4564 896
rect 1540 840 2604 868
rect 3500 840 4536 868
rect 1596 812 2744 840
rect 3332 812 4508 840
rect 1624 784 4452 812
rect 1652 756 4424 784
rect 1708 728 4368 756
rect 1764 700 4340 728
rect 1792 672 4284 700
rect 1848 644 4228 672
rect 1904 616 4172 644
rect 1960 588 4144 616
rect 2016 560 4060 588
rect 2072 532 4004 560
rect 2128 504 3948 532
rect 2212 476 3864 504
rect 2296 448 3780 476
rect 2380 420 3696 448
rect 2492 392 3584 420
rect 2632 364 3444 392
<< end >>
