magic
tech sky130A
magscale 1 2
timestamp 1711565985
<< error_p >>
rect 19863 24036 19909 24048
rect 19863 23998 19869 24036
rect 19863 23986 19909 23998
rect 19863 23908 19909 23920
rect 19863 23870 19869 23908
rect 19863 23858 19909 23870
rect 19863 23780 19909 23792
rect 19863 23742 19869 23780
rect 19863 23730 19909 23742
rect 19863 23652 19909 23664
rect 19863 23614 19869 23652
rect 19863 23602 19909 23614
rect 19863 23524 19909 23536
rect 19863 23486 19869 23524
rect 19863 23474 19909 23486
rect 19863 23396 19909 23408
rect 19863 23358 19869 23396
rect 19863 23346 19909 23358
rect 19863 23268 19909 23280
rect 19863 23230 19869 23268
rect 19863 23218 19909 23230
rect 19863 23140 19909 23152
rect 19863 23102 19869 23140
rect 19863 23090 19909 23102
rect 30173 22164 30219 22176
rect 32301 22164 32347 22176
rect 32409 22164 32455 22176
rect 34537 22164 34583 22176
rect 34645 22164 34691 22176
rect 36773 22164 36819 22176
rect 30173 22126 30179 22164
rect 32301 22126 32307 22164
rect 32409 22126 32415 22164
rect 34537 22126 34543 22164
rect 34645 22126 34651 22164
rect 36773 22126 36779 22164
rect 30173 22114 30219 22126
rect 32301 22114 32347 22126
rect 32409 22114 32455 22126
rect 34537 22114 34583 22126
rect 34645 22114 34691 22126
rect 36773 22114 36819 22126
rect 32569 20606 32615 20618
rect 32677 20606 32723 20618
rect 34805 20606 34851 20618
rect 34913 20606 34959 20618
rect 37041 20606 37087 20618
rect 32569 20568 32575 20606
rect 32677 20568 32683 20606
rect 34805 20568 34811 20606
rect 34913 20568 34919 20606
rect 37041 20568 37047 20606
rect 32569 20556 32615 20568
rect 32677 20556 32723 20568
rect 34805 20556 34851 20568
rect 34913 20556 34959 20568
rect 37041 20556 37087 20568
rect 11400 19292 11446 19304
rect 11928 19292 11974 19304
rect 11400 19258 11406 19292
rect 11928 19258 11934 19292
rect 11400 19246 11446 19258
rect 11928 19246 11974 19258
rect 11400 18976 11446 18988
rect 11928 18976 11974 18988
rect 11400 18942 11406 18976
rect 11928 18942 11934 18976
rect 11400 18930 11446 18942
rect 11928 18930 11974 18942
rect 11500 18518 11546 18530
rect 11810 18518 11856 18530
rect 11500 18484 11506 18518
rect 11810 18484 11816 18518
rect 11500 18472 11546 18484
rect 11810 18472 11856 18484
rect 11500 18202 11546 18214
rect 11810 18202 11856 18214
rect 11500 18168 11506 18202
rect 11810 18168 11816 18202
rect 11500 18156 11546 18168
rect 11810 18156 11856 18168
rect 4726 14974 4772 14986
rect 5254 14974 5300 14986
rect 4726 14940 4732 14974
rect 5254 14940 5260 14974
rect 4726 14928 4772 14940
rect 5254 14928 5300 14940
rect 4726 14658 4772 14670
rect 5254 14658 5300 14670
rect 4726 14624 4732 14658
rect 5254 14624 5260 14658
rect 4726 14612 4772 14624
rect 5254 14612 5300 14624
rect 4826 14200 4872 14212
rect 5136 14200 5182 14212
rect 4826 14166 4832 14200
rect 5136 14166 5142 14200
rect 4826 14154 4872 14166
rect 5136 14154 5182 14166
rect 4826 13884 4872 13896
rect 5136 13884 5182 13896
rect 4826 13850 4832 13884
rect 5136 13850 5142 13884
rect 4826 13838 4872 13850
rect 5136 13838 5182 13850
rect 24246 4892 24308 4898
rect 24246 4858 24258 4892
rect 24246 4852 24308 4858
rect 24246 3782 24308 3788
rect 24246 3748 24258 3782
rect 24246 3742 24308 3748
rect 24246 3674 24308 3680
rect 24246 3640 24258 3674
rect 24246 3634 24308 3640
rect 24246 2564 24308 2570
rect 24246 2530 24258 2564
rect 24246 2524 24308 2530
rect 24246 2456 24308 2462
rect 24246 2422 24258 2456
rect 24246 2416 24308 2422
rect 24246 1346 24308 1352
rect 24246 1312 24258 1346
rect 24246 1306 24308 1312
rect 24246 1238 24308 1244
rect 24246 1204 24258 1238
rect 24246 1198 24308 1204
rect 24246 128 24308 134
rect 24246 94 24258 128
rect 24246 88 24308 94
<< error_s >>
rect 8493 3459 8714 3469
rect 8747 2831 8968 3459
rect 9148 2421 9169 3227
rect 9176 2821 9423 3459
rect 9176 2393 9197 2821
rect 9577 2421 9598 3227
rect 9605 2821 9852 3459
rect 9605 2393 9626 2821
rect 10006 2421 10027 3227
rect 10034 2821 10281 3459
rect 10034 2393 10055 2821
rect 10435 2421 10456 3227
rect 10463 2821 10710 3459
rect 10463 2393 10484 2821
rect 10864 2421 10885 3227
rect 10892 2821 11139 3459
rect 10892 2393 10913 2821
rect 17565 1811 17599 1829
rect 17529 352 17599 1811
rect 17529 347 17600 352
rect 17529 311 17582 347
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use comp_n  X_COMP_N
timestamp 1711057506
transform -1 0 71974 0 1 4920
box 18500 1578 24043 5238
use comp_p  X_COMP_P1
timestamp 1711565985
transform 1 0 26493 0 1 18384
box -3598 1576 2410 5166
use inv  X_INV1
timestamp 1711045747
transform 1 0 8352 0 1 1649
box -60 547 369 1820
use inv  X_INV2[0]
timestamp 1711045747
transform 1 0 9236 0 1 1639
box -60 547 369 1820
use inv  X_INV2[1]
timestamp 1711045747
transform 1 0 8807 0 1 1639
box -60 547 369 1820
use inv  X_INV3[0]
timestamp 1711045747
transform 1 0 10952 0 1 1639
box -60 547 369 1820
use inv  X_INV3[1]
timestamp 1711045747
transform 1 0 10523 0 1 1639
box -60 547 369 1820
use inv  X_INV3[2]
timestamp 1711045747
transform 1 0 10094 0 1 1639
box -60 547 369 1820
use inv  X_INV3[3]
timestamp 1711045747
transform 1 0 9665 0 1 1639
box -60 547 369 1820
use sr_latch  X_SR_LATCH
timestamp 1711045747
transform 1 0 8745 0 1 14056
box -4457 -2000 3703 5706
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_bias
timestamp 1711041810
transform 1 0 17286 0 1 1045
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_44Y62X  XMn_discharge
timestamp 1711041017
transform 1 0 24277 0 1 2493
box -231 -2537 2431 2537
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_bias
timestamp 1711036998
transform 1 0 17825 0 1 1501
box -296 -1219 296 1219
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_1
timestamp 1711037431
transform 1 0 10561 0 1 -2770
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_2
timestamp 1711037431
transform 1 0 13413 0 1 -2446
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_3
timestamp 1711037431
transform 1 0 14119 0 1 -2418
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_4
timestamp 1711037431
transform 1 0 14973 0 1 -2418
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bot
timestamp 1711037431
transform 1 0 9795 0 1 -2828
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_mid
timestamp 1711037431
transform 1 0 9089 0 1 -2946
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_top
timestamp 1711037431
transform 1 0 8383 0 1 -2976
box -307 -1282 307 1282
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 DO_OUT
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 V_DISCH_O
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 V_THRESH_I
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 V_TRIG_B_I
port 5 nsew
<< end >>
