magic
tech sky130A
magscale 1 2
timestamp 1711745511
<< nwell >>
rect 20680 18281 23158 18315
<< pwell >>
rect 20680 17271 23166 17305
<< psubdiff >>
rect 20680 17271 23166 17305
<< nsubdiff >>
rect 24103 19828 28001 19886
rect 20680 18281 23158 18315
<< locali >>
rect 21942 23276 22918 23410
rect 21852 22844 23008 22938
rect 20679 17190 23156 17305
rect 20679 17156 20810 17190
rect 22966 17156 23156 17190
<< viali >>
rect 20810 17156 22966 17190
rect 20696 16384 20748 17094
<< metal1 >>
rect 20631 23478 20641 23878
rect 28516 23478 28587 23878
rect 21942 23472 22918 23478
rect 22056 23276 22804 23472
rect 22962 23062 23030 23080
rect 20798 21930 21230 22720
rect 22598 22438 23030 23062
rect 23246 22282 23322 22288
rect 23246 22224 23252 22282
rect 23316 22279 23322 22282
rect 23316 22227 23498 22279
rect 23316 22224 23322 22227
rect 23246 22218 23322 22224
rect 20798 20914 21230 21704
rect 22598 21422 23030 22212
rect 22598 20514 23030 21196
rect 25275 20548 25285 20604
rect 25661 20548 25671 20604
rect 26475 20548 26485 20604
rect 26861 20548 26871 20604
rect 22938 20368 23030 20514
rect 23352 20372 23428 20378
rect 23352 20368 23358 20372
rect 22938 20316 23358 20368
rect 22938 20304 23030 20316
rect 23352 20314 23358 20316
rect 23422 20314 23428 20372
rect 23352 20308 23428 20314
rect 20909 20196 22885 20288
rect 20800 20140 20810 20196
rect 22984 20140 22994 20196
rect 26219 19916 26229 20030
rect 20798 19510 21230 19862
rect 22598 19688 22608 19876
rect 23018 19688 23028 19876
rect 23522 19798 26229 19916
rect 26219 19685 26229 19798
rect 26790 19916 26800 20030
rect 26790 19798 28576 19916
rect 26790 19685 26800 19798
rect 23246 19512 23322 19518
rect 23246 19510 23252 19512
rect 20798 19458 23252 19510
rect 20798 19100 21230 19458
rect 23246 19454 23252 19458
rect 23316 19454 23322 19512
rect 23246 19448 23322 19454
rect 20272 18590 21230 18872
rect 22598 18646 23030 19352
rect 25275 19110 25285 19166
rect 25661 19110 25671 19166
rect 26475 19110 26485 19166
rect 26861 19110 26871 19166
rect 23246 18650 23322 18656
rect 23246 18646 23252 18650
rect 22598 18594 23252 18646
rect 22598 18590 23030 18594
rect 23246 18592 23252 18594
rect 23316 18592 23322 18650
rect 20272 17305 20554 18590
rect 23246 18586 23322 18592
rect 24432 18538 24442 18590
rect 25395 18538 25405 18590
rect 20646 18281 20656 18333
rect 23181 18281 23191 18333
rect 23246 17490 23322 17496
rect 23246 17432 23252 17490
rect 23316 17488 23322 17490
rect 23316 17436 23490 17488
rect 23316 17432 23322 17436
rect 23246 17426 23322 17432
rect 20272 17271 23166 17305
rect 20272 17190 23156 17271
rect 20272 17156 20810 17190
rect 22966 17156 23156 17190
rect 20272 15831 20554 17156
rect 20667 17106 20748 17156
rect 20798 17150 22978 17156
rect 20667 17094 20754 17106
rect 20667 16384 20696 17094
rect 20748 16384 20754 17094
rect 20810 16448 20856 17030
rect 22920 16448 22966 17030
rect 20667 16372 20754 16384
rect 20667 16338 20748 16372
rect 20667 16276 28610 16338
rect 20667 16236 28614 16276
rect 20667 15836 20677 16236
rect 28613 15836 28623 16236
<< via1 >>
rect 20641 23478 28516 23878
rect 23252 22224 23316 22282
rect 25285 20548 25661 20604
rect 26485 20548 26861 20604
rect 23358 20314 23422 20372
rect 20810 20140 22984 20196
rect 22608 19688 23018 19876
rect 26229 19685 26790 20030
rect 23252 19454 23316 19512
rect 25285 19110 25661 19166
rect 26485 19110 26861 19166
rect 23252 18592 23316 18650
rect 24442 18538 25395 18590
rect 20656 18281 23181 18333
rect 23252 17432 23316 17490
rect 20677 15836 28613 16236
<< metal2 >>
rect 20641 23878 28577 23888
rect 28516 23478 28578 23878
rect 20641 23468 28577 23478
rect 23246 22282 23322 22288
rect 23246 22224 23252 22282
rect 23316 22224 23322 22282
rect 23246 22218 23322 22224
rect 20810 20196 22984 20206
rect 20810 20130 22984 20140
rect 22608 19876 23018 19886
rect 22608 19678 23018 19688
rect 23258 19518 23310 22218
rect 25285 20604 25661 20614
rect 25285 20538 25661 20548
rect 26485 20604 26861 20614
rect 26485 20538 26861 20548
rect 23352 20372 23428 20378
rect 23352 20314 23358 20372
rect 23422 20314 23428 20372
rect 23352 20308 23428 20314
rect 23364 19984 23416 20308
rect 26229 20030 26790 20040
rect 23364 19932 23492 19984
rect 23364 19782 23416 19932
rect 23364 19730 23490 19782
rect 26229 19675 26790 19685
rect 23246 19512 23322 19518
rect 23246 19454 23252 19512
rect 23316 19454 23322 19512
rect 23246 19448 23322 19454
rect 25276 19166 25670 19174
rect 25276 19110 25285 19166
rect 25661 19110 25670 19166
rect 25276 19100 25670 19110
rect 26476 19166 26870 19174
rect 26476 19110 26485 19166
rect 26861 19110 26870 19166
rect 26476 19100 26870 19110
rect 23246 18650 23322 18656
rect 23246 18592 23252 18650
rect 23316 18592 23322 18650
rect 23246 18586 23322 18592
rect 24442 18594 25395 18604
rect 20656 18337 23181 18347
rect 20656 18271 23181 18281
rect 23258 17496 23310 18586
rect 24442 18528 25395 18538
rect 23246 17490 23322 17496
rect 23246 17432 23252 17490
rect 23316 17432 23322 17490
rect 23246 17426 23322 17432
rect 20677 16236 28613 16246
rect 20677 15826 28613 15836
<< via2 >>
rect 20641 23478 28166 23878
rect 20810 20140 22984 20196
rect 22608 19688 23018 19876
rect 25285 20548 25661 20604
rect 26485 20548 26861 20604
rect 26229 19685 26790 20030
rect 25285 19110 25661 19166
rect 26485 19110 26861 19166
rect 24442 18590 25395 18594
rect 20656 18333 23181 18337
rect 20656 18281 23181 18333
rect 24442 18538 25395 18590
rect 20677 15836 28166 16236
<< metal3 >>
rect 20631 23878 28613 23883
rect 20631 23874 20641 23878
rect 20428 23478 20641 23874
rect 28166 23478 28613 23878
rect 20428 23474 28613 23478
rect 20631 23473 28613 23474
rect 20428 21123 26861 21523
rect 25285 20609 25661 21123
rect 26485 20609 26861 21123
rect 25275 20604 25671 20609
rect 25275 20548 25285 20604
rect 25661 20548 25671 20604
rect 25275 20543 25671 20548
rect 26475 20604 26871 20609
rect 26475 20548 26485 20604
rect 26861 20548 26871 20604
rect 26475 20543 26871 20548
rect 20800 20196 22994 20201
rect 20800 20140 20810 20196
rect 22984 20140 22994 20196
rect 20800 20068 22994 20140
rect 25285 20068 25661 20543
rect 26485 20120 26861 20543
rect 26485 20068 26860 20120
rect 20428 20030 26860 20068
rect 20428 19876 26229 20030
rect 20428 19688 22608 19876
rect 23018 19688 26229 19876
rect 20428 19685 26229 19688
rect 26790 19685 26860 20030
rect 20428 19650 26860 19685
rect 20428 19648 26861 19650
rect 25285 19171 25661 19648
rect 26485 19171 26861 19648
rect 25275 19166 25671 19171
rect 25275 19110 25285 19166
rect 25661 19110 25671 19166
rect 25275 19105 25671 19110
rect 26475 19166 26871 19171
rect 26475 19110 26485 19166
rect 26861 19110 26871 19166
rect 26475 19105 26871 19110
rect 25285 18599 25661 19105
rect 24432 18594 25661 18599
rect 24432 18592 24442 18594
rect 20428 18538 24442 18592
rect 25395 18592 25661 18594
rect 26485 18630 26861 19105
rect 26485 18592 26860 18630
rect 25395 18538 26860 18592
rect 20428 18337 26860 18538
rect 20428 18281 20656 18337
rect 23181 18281 26860 18337
rect 20428 18192 26860 18281
rect 28213 16241 28613 23473
rect 20667 16236 28613 16241
rect 20667 16231 20677 16236
rect 20428 15836 20677 16231
rect 28166 15894 28613 16236
rect 28166 15836 28623 15894
rect 20428 15831 28623 15836
use comp_p  X_COMP_P_BOTTOM
timestamp 1711732688
transform 1 0 26492 0 1 14702
box -3002 1462 2120 5166
use comp_p  X_COMP_P_TOP
timestamp 1711732688
transform 1 0 26493 0 -1 25012
box -3002 1462 2120 5166
use inv  X_INV1
timestamp 1711732688
transform 1 0 20381 0 1 16477
box 978 788 1260 1874
use inv  X_INV2[0]
timestamp 1711732688
transform 1 0 20906 0 1 16477
box 978 788 1260 1874
use inv  X_INV2[1]
timestamp 1711732688
transform 1 0 20643 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[0]
timestamp 1711732688
transform 1 0 21958 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[1]
timestamp 1711732688
transform 1 0 21695 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[2]
timestamp 1711732688
transform 1 0 21432 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[3]
timestamp 1711732688
transform 1 0 21169 0 1 16477
box 978 788 1260 1874
use sr_latch  X_SR_LATCH
timestamp 1711732688
transform -1 0 15343 0 1 16911
box -6020 354 -5267 1440
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_bias
timestamp 1711732688
transform 0 1 22430 -1 0 23164
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_NVJ7JE  XMn_discharge
timestamp 1711736161
transform 0 1 21888 -1 0 16739
box -487 -1210 487 1210
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_bias
timestamp 1711732688
transform 0 1 21897 -1 0 20400
box -296 -1219 296 1219
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_1
timestamp 1711732688
transform 0 1 21914 1 0 21055
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_2
timestamp 1711732688
transform 0 1 21914 1 0 21563
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_3
timestamp 1711732688
transform 0 1 21914 1 0 22071
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_4
timestamp 1711732688
transform 0 1 21914 1 0 22579
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bot
timestamp 1711732688
transform 0 1 21914 -1 0 18731
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_mid
timestamp 1711732688
transform 0 1 21914 -1 0 19239
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_top
timestamp 1711732688
transform 0 1 21914 -1 0 19747
box -307 -1282 307 1282
<< end >>
