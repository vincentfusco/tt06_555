magic
tech sky130A
magscale 1 2
timestamp 1711658383
<< nwell >>
rect -3002 4716 2120 5166
rect -3002 4710 -566 4716
rect -518 4710 2120 4716
rect -3002 2542 2120 4710
<< pwell >>
rect -3002 1464 2120 2542
<< pmoslvt >>
rect -2577 3672 -578 3742
rect -2577 3432 -578 3502
rect -2577 3192 -578 3262
rect -2577 2952 -578 3022
rect -305 3672 1694 3742
rect -305 3432 1694 3502
rect -305 3192 1694 3262
rect -305 2952 1694 3022
<< pdiff >>
rect -2577 3788 -578 3800
rect -2577 3754 -2565 3788
rect -590 3754 -578 3788
rect -2577 3742 -578 3754
rect -2577 3660 -578 3672
rect -2577 3626 -2565 3660
rect -590 3626 -578 3660
rect -2577 3614 -578 3626
rect -2577 3548 -578 3560
rect -2577 3514 -2565 3548
rect -590 3514 -578 3548
rect -2577 3502 -578 3514
rect -2577 3420 -578 3432
rect -2577 3386 -2565 3420
rect -590 3386 -578 3420
rect -2577 3374 -578 3386
rect -2577 3308 -578 3320
rect -2577 3274 -2565 3308
rect -590 3274 -578 3308
rect -2577 3262 -578 3274
rect -2577 3180 -578 3192
rect -2577 3146 -2565 3180
rect -590 3146 -578 3180
rect -2577 3134 -578 3146
rect -2577 3068 -578 3080
rect -2577 3034 -2565 3068
rect -590 3034 -578 3068
rect -2577 3022 -578 3034
rect -2577 2940 -578 2952
rect -2577 2906 -2565 2940
rect -590 2906 -578 2940
rect -2577 2894 -578 2906
rect -305 3788 1694 3800
rect -305 3754 -293 3788
rect 1682 3754 1694 3788
rect -305 3742 1694 3754
rect -305 3660 1694 3672
rect -305 3626 -293 3660
rect 1686 3626 1694 3660
rect -305 3614 1694 3626
rect -305 3548 1694 3560
rect -305 3514 -293 3548
rect 1682 3514 1694 3548
rect -305 3502 1694 3514
rect -305 3420 1694 3432
rect -305 3386 -293 3420
rect 1682 3386 1694 3420
rect -305 3374 1694 3386
rect -305 3308 1694 3320
rect -305 3274 -293 3308
rect 1682 3274 1694 3308
rect -305 3262 1694 3274
rect -305 3180 1694 3192
rect -305 3146 -293 3180
rect 1686 3146 1694 3180
rect -305 3134 1694 3146
rect -305 3068 1694 3080
rect -305 3034 -293 3068
rect 1682 3034 1694 3068
rect -305 3022 1694 3034
rect -305 2940 1694 2952
rect -305 2906 -293 2940
rect 1682 2906 1694 2940
rect -305 2894 1694 2906
<< pdiffc >>
rect -2565 3754 -590 3788
rect -2565 3626 -590 3660
rect -2565 3514 -590 3548
rect -2565 3386 -590 3420
rect -2565 3274 -590 3308
rect -2565 3146 -590 3180
rect -2565 3034 -590 3068
rect -2565 2906 -590 2940
rect -293 3754 1682 3788
rect -293 3626 1686 3660
rect -293 3514 1682 3548
rect -293 3386 1682 3420
rect -293 3274 1682 3308
rect -293 3146 1686 3180
rect -293 3034 1682 3068
rect -293 2906 1682 2940
<< nsubdiff >>
rect -2730 3854 -2650 3888
rect -497 3854 -378 3888
rect 1775 3854 1847 3888
rect -2730 3792 -2696 3854
rect -458 3792 -424 3854
rect -2730 2840 -2696 2902
rect 1813 3792 1847 3854
rect -458 2840 -424 2902
rect 1813 2840 1847 2902
rect -2730 2806 -2650 2840
rect -497 2806 -378 2840
rect 1775 2806 1847 2840
<< nsubdiffcont >>
rect -2650 3854 -497 3888
rect -378 3854 1775 3888
rect -2730 2902 -2696 3792
rect -458 2902 -424 3792
rect 1813 2902 1847 3792
rect -2650 2806 -497 2840
rect -378 2806 1775 2840
<< poly >>
rect -2674 3726 -2577 3742
rect -2674 3688 -2658 3726
rect -2624 3688 -2577 3726
rect -2674 3672 -2577 3688
rect -578 3726 -481 3742
rect -578 3688 -531 3726
rect -497 3688 -481 3726
rect -578 3672 -481 3688
rect -2674 3486 -2577 3502
rect -2674 3448 -2658 3486
rect -2624 3448 -2577 3486
rect -2674 3432 -2577 3448
rect -578 3486 -481 3502
rect -578 3448 -531 3486
rect -497 3448 -481 3486
rect -578 3432 -481 3448
rect -2674 3246 -2577 3262
rect -2674 3208 -2658 3246
rect -2624 3208 -2577 3246
rect -2674 3192 -2577 3208
rect -578 3246 -481 3262
rect -578 3208 -531 3246
rect -497 3208 -481 3246
rect -578 3192 -481 3208
rect -2674 3006 -2577 3022
rect -2674 2968 -2658 3006
rect -2624 2968 -2577 3006
rect -2674 2952 -2577 2968
rect -578 3006 -481 3022
rect -578 2968 -531 3006
rect -497 2968 -481 3006
rect -578 2952 -481 2968
rect -402 3726 -305 3742
rect -402 3688 -386 3726
rect -352 3688 -305 3726
rect -402 3672 -305 3688
rect 1694 3726 1791 3742
rect 1694 3688 1741 3726
rect 1775 3688 1791 3726
rect 1694 3672 1791 3688
rect -402 3486 -305 3502
rect -402 3448 -386 3486
rect -352 3448 -305 3486
rect -402 3432 -305 3448
rect 1694 3486 1791 3502
rect 1694 3448 1741 3486
rect 1775 3448 1791 3486
rect 1694 3432 1791 3448
rect -402 3246 -305 3262
rect -402 3208 -386 3246
rect -352 3208 -305 3246
rect -402 3192 -305 3208
rect 1694 3246 1791 3262
rect 1694 3208 1741 3246
rect 1775 3208 1791 3246
rect 1694 3192 1791 3208
rect -402 3006 -305 3022
rect -402 2968 -386 3006
rect -352 2968 -305 3006
rect -402 2952 -305 2968
rect 1694 3006 1791 3022
rect 1694 2968 1741 3006
rect 1775 2968 1791 3006
rect 1694 2952 1791 2968
<< polycont >>
rect -2658 3688 -2624 3726
rect -531 3688 -497 3726
rect -2658 3448 -2624 3486
rect -531 3448 -497 3486
rect -2658 3208 -2624 3246
rect -531 3208 -497 3246
rect -2658 2968 -2624 3006
rect -531 2968 -497 3006
rect -386 3688 -352 3726
rect 1741 3688 1775 3726
rect -386 3448 -352 3486
rect 1741 3448 1775 3486
rect -386 3208 -352 3246
rect 1741 3208 1775 3246
rect -386 2968 -352 3006
rect 1741 2968 1775 3006
<< locali >>
rect -2968 4644 -2354 5096
rect 1474 4646 2084 5096
rect 728 4644 2084 4646
rect -2968 4522 2084 4644
rect -2968 4070 -1568 4522
rect -1407 4408 569 4522
rect 728 4070 2084 4522
rect -2968 3888 2084 4070
rect -2968 3854 -2650 3888
rect -497 3854 -378 3888
rect 1775 3854 2084 3888
rect -2968 3792 -2696 3854
rect -2968 2902 -2730 3792
rect -458 3792 -424 3854
rect -2581 3754 -2565 3788
rect -590 3754 -574 3788
rect -2658 3726 -2624 3742
rect -2658 3672 -2624 3688
rect -531 3726 -497 3742
rect -531 3672 -497 3688
rect -2581 3626 -2565 3660
rect -590 3626 -574 3660
rect -2581 3514 -2565 3548
rect -590 3514 -574 3548
rect -2658 3486 -2624 3502
rect -2658 3432 -2624 3448
rect -531 3486 -497 3502
rect -531 3432 -497 3448
rect -2581 3386 -2565 3420
rect -590 3386 -574 3420
rect -2581 3274 -2565 3308
rect -590 3274 -574 3308
rect -2658 3246 -2624 3262
rect -2658 3192 -2624 3208
rect -531 3246 -497 3262
rect -531 3192 -497 3208
rect -2581 3146 -2565 3180
rect -590 3146 -574 3180
rect -2581 3034 -2565 3068
rect -590 3034 -574 3068
rect -2658 3006 -2624 3022
rect -2658 2952 -2624 2968
rect -531 3006 -497 3022
rect -531 2952 -497 2968
rect -2581 2906 -2565 2940
rect -590 2906 -574 2940
rect -2968 2840 -2696 2902
rect 1813 3792 2084 3854
rect -309 3754 -293 3788
rect 1682 3754 1698 3788
rect -386 3726 -352 3742
rect -386 3672 -352 3688
rect 1741 3726 1775 3742
rect 1546 3660 1690 3676
rect 1741 3672 1775 3688
rect -309 3626 -293 3660
rect 1686 3626 1698 3660
rect 1546 3608 1690 3626
rect -309 3514 -293 3548
rect 1682 3514 1698 3548
rect -386 3486 -352 3502
rect -386 3432 -352 3448
rect 1741 3486 1775 3502
rect 1741 3432 1775 3448
rect -309 3386 -293 3420
rect 1682 3386 1698 3420
rect -309 3274 -293 3308
rect 1682 3274 1698 3308
rect -386 3246 -352 3262
rect -386 3192 -352 3208
rect 1741 3246 1775 3262
rect 1546 3180 1690 3196
rect 1741 3192 1775 3208
rect -309 3146 -293 3180
rect 1686 3146 1698 3180
rect 1546 3128 1690 3146
rect -309 3034 -293 3068
rect 1682 3034 1698 3068
rect -386 3006 -352 3022
rect -386 2952 -352 2968
rect 1741 3006 1775 3022
rect 1741 2952 1775 2968
rect -309 2906 -293 2940
rect 1682 2906 1698 2940
rect -458 2840 -424 2902
rect 1847 2902 2084 3792
rect 1813 2840 2084 2902
rect -2968 2806 -2650 2840
rect -497 2806 -378 2840
rect 1775 2806 2084 2840
rect -2780 2102 -2004 2140
rect -1610 2102 -634 2134
rect -216 2102 760 2134
rect 1122 2102 1898 2140
rect -2968 1986 2084 2102
rect -2968 1534 -1818 1986
rect 936 1534 2084 1986
<< viali >>
rect -2968 5096 2084 5130
rect -2565 3754 -590 3788
rect -2658 3688 -2624 3726
rect -531 3688 -497 3726
rect -2565 3626 -590 3660
rect -2565 3514 -590 3548
rect -2658 3448 -2624 3486
rect -531 3448 -497 3486
rect -2565 3386 -590 3420
rect -2565 3274 -590 3308
rect -2658 3208 -2624 3246
rect -531 3208 -497 3246
rect -2565 3146 -590 3180
rect -2565 3034 -590 3068
rect -2658 2968 -2624 3006
rect -531 2968 -497 3006
rect -2565 2906 -590 2940
rect -293 3754 1682 3788
rect -386 3688 -352 3726
rect 1741 3688 1775 3726
rect -293 3626 1686 3660
rect -293 3514 1682 3548
rect -386 3448 -352 3486
rect 1741 3448 1775 3486
rect -293 3386 1682 3420
rect -293 3274 1682 3308
rect -386 3208 -352 3246
rect 1741 3208 1775 3246
rect -293 3146 1686 3180
rect -293 3034 1682 3068
rect -386 2968 -352 3006
rect 1741 2968 1775 3006
rect -293 2906 1682 2940
rect -2968 1500 2084 1534
<< metal1 >>
rect -3002 5130 2120 5166
rect -3002 5096 -2968 5130
rect 2084 5096 2120 5130
rect -3002 5090 2120 5096
rect -3002 4644 -2354 5090
rect -2195 4982 -619 5090
rect -263 4982 1313 5090
rect -566 4954 -520 4966
rect -566 4898 -322 4954
rect -2252 4846 1406 4898
rect -566 4786 -322 4846
rect -2294 4768 -2248 4780
rect -566 4768 -520 4786
rect -2294 4716 -2196 4768
rect -620 4716 -520 4768
rect -274 4716 -264 4768
rect 1312 4716 1322 4768
rect 1472 4644 2120 5090
rect -3002 4572 2120 4644
rect -1520 4212 -1510 4380
rect -1458 4212 -1448 4380
rect 608 4212 618 4380
rect 670 4212 680 4380
rect -1417 4144 -1407 4196
rect 569 4144 579 4196
rect -3002 3924 -2666 3976
rect -2614 3924 -540 3976
rect -488 3924 1858 3976
rect -720 3796 -576 3802
rect -720 3794 -712 3796
rect -2577 3788 -712 3794
rect -2577 3754 -2565 3788
rect -2577 3748 -712 3754
rect -720 3744 -712 3748
rect -586 3744 -576 3796
rect -304 3794 -296 3796
rect -305 3748 -296 3794
rect -170 3794 -164 3796
rect -170 3788 1694 3794
rect 1682 3754 1694 3788
rect -720 3738 -576 3744
rect -304 3744 -296 3748
rect -170 3748 1694 3754
rect -170 3744 -86 3748
rect -304 3742 -86 3744
rect -2668 3726 -2612 3738
rect -2738 3688 -2658 3726
rect -2624 3688 -2612 3726
rect -2738 3246 -2700 3688
rect -2668 3676 -2612 3688
rect -540 3726 -486 3738
rect -540 3688 -531 3726
rect -497 3688 -486 3726
rect -540 3676 -486 3688
rect -396 3726 -340 3738
rect -396 3688 -386 3726
rect -352 3688 -340 3726
rect -396 3676 -340 3688
rect 1732 3726 1786 3738
rect 1820 3726 1858 3924
rect 1732 3688 1741 3726
rect 1775 3688 1858 3726
rect 1732 3676 1786 3688
rect -2572 3668 -2428 3674
rect 1546 3668 1690 3676
rect -2572 3666 -2564 3668
rect -2577 3660 -2564 3666
rect -2438 3666 -2428 3668
rect -306 3666 -86 3668
rect 1546 3666 1556 3668
rect -2438 3660 -578 3666
rect -2577 3626 -2565 3660
rect -590 3626 -578 3660
rect -2577 3620 -2564 3626
rect -2572 3616 -2564 3620
rect -2438 3620 -578 3626
rect -306 3660 1556 3666
rect 1682 3666 1690 3668
rect 1682 3660 1694 3666
rect -306 3626 -293 3660
rect 1686 3626 1694 3660
rect -306 3620 1556 3626
rect -2438 3616 -2428 3620
rect -306 3616 -86 3620
rect 1546 3616 1556 3620
rect 1682 3620 1694 3626
rect 1682 3616 1690 3620
rect -2572 3610 -2428 3616
rect 1546 3608 1690 3616
rect -720 3556 -576 3562
rect -720 3554 -712 3556
rect -2577 3548 -712 3554
rect -2577 3514 -2565 3548
rect -2577 3508 -712 3514
rect -720 3504 -712 3508
rect -586 3504 -576 3556
rect -304 3556 -160 3564
rect -304 3554 -296 3556
rect -305 3508 -296 3554
rect -170 3554 -160 3556
rect -170 3548 1694 3554
rect 1682 3514 1694 3548
rect -720 3498 -576 3504
rect -304 3504 -296 3508
rect -170 3508 1694 3514
rect -170 3504 -160 3508
rect -2672 3494 -2608 3498
rect -2672 3442 -2666 3494
rect -2614 3442 -2608 3494
rect -2672 3436 -2608 3442
rect -548 3492 -480 3502
rect -548 3440 -540 3492
rect -488 3440 -480 3492
rect -548 3432 -480 3440
rect -402 3492 -334 3502
rect -304 3498 -160 3504
rect -402 3440 -392 3492
rect -340 3440 -334 3492
rect -402 3432 -334 3440
rect 1726 3494 1792 3504
rect 1726 3442 1732 3494
rect 1784 3442 1792 3494
rect 1726 3432 1792 3442
rect -2332 3428 -2188 3432
rect -2332 3426 -2324 3428
rect -2577 3420 -2324 3426
rect -2198 3426 -2188 3428
rect 1306 3426 1316 3428
rect -2198 3420 -578 3426
rect -2577 3386 -2565 3420
rect -590 3386 -578 3420
rect -2577 3380 -2324 3386
rect -2332 3376 -2324 3380
rect -2198 3380 -578 3386
rect -305 3420 1316 3426
rect 1442 3426 1450 3428
rect 1442 3420 1694 3426
rect -305 3386 -293 3420
rect 1682 3386 1694 3420
rect -305 3380 1316 3386
rect -2198 3376 -2188 3380
rect 1306 3376 1316 3380
rect 1442 3380 1694 3386
rect 1442 3376 1450 3380
rect -2332 3370 -2188 3376
rect -720 3316 -576 3322
rect -720 3314 -712 3316
rect -2577 3308 -712 3314
rect -2577 3274 -2565 3308
rect -2577 3268 -712 3274
rect -720 3264 -712 3268
rect -586 3264 -576 3316
rect -304 3316 -160 3324
rect -304 3314 -296 3316
rect -305 3268 -296 3314
rect -170 3314 -160 3316
rect -170 3308 1694 3314
rect 1682 3274 1694 3308
rect -720 3258 -576 3264
rect -304 3264 -296 3268
rect -170 3268 1694 3274
rect -170 3264 -94 3268
rect -304 3262 -94 3264
rect -2668 3246 -2612 3258
rect -2738 3208 -2658 3246
rect -2624 3208 -2612 3246
rect -2738 2786 -2700 3208
rect -2668 3196 -2612 3208
rect -540 3246 -486 3258
rect -540 3208 -531 3246
rect -497 3208 -486 3246
rect -540 3196 -486 3208
rect -396 3246 -340 3258
rect -396 3208 -386 3246
rect -352 3208 -340 3246
rect -396 3196 -340 3208
rect 1732 3246 1786 3258
rect 1820 3246 1858 3688
rect 1732 3208 1741 3246
rect 1775 3208 1858 3246
rect 1732 3196 1786 3208
rect -2572 3188 -2428 3194
rect 1546 3188 1690 3196
rect -2572 3186 -2564 3188
rect -2577 3180 -2564 3186
rect -2438 3186 -2428 3188
rect -306 3186 -94 3188
rect 1546 3186 1556 3188
rect -2438 3180 -578 3186
rect -2577 3146 -2565 3180
rect -590 3146 -578 3180
rect -2577 3140 -2564 3146
rect -2572 3136 -2564 3140
rect -2438 3140 -578 3146
rect -306 3180 1556 3186
rect 1682 3186 1690 3188
rect 1682 3180 1694 3186
rect -306 3146 -293 3180
rect 1686 3146 1694 3180
rect -306 3140 1556 3146
rect -2438 3136 -2428 3140
rect -306 3136 -94 3140
rect 1546 3136 1556 3140
rect 1682 3140 1694 3146
rect 1682 3136 1690 3140
rect -2572 3130 -2428 3136
rect 1546 3128 1690 3136
rect -720 3076 -576 3082
rect -720 3074 -712 3076
rect -2577 3068 -712 3074
rect -2577 3034 -2565 3068
rect -2577 3028 -712 3034
rect -720 3024 -712 3028
rect -586 3024 -576 3076
rect -304 3076 -160 3084
rect -304 3074 -296 3076
rect -305 3028 -296 3074
rect -170 3074 -160 3076
rect -170 3068 1694 3074
rect 1682 3034 1694 3068
rect -720 3018 -576 3024
rect -304 3024 -296 3028
rect -170 3028 1694 3034
rect -170 3024 -160 3028
rect -2672 3014 -2608 3018
rect -2672 2962 -2666 3014
rect -2614 2962 -2608 3014
rect -2672 2956 -2608 2962
rect -548 3012 -480 3022
rect -548 2960 -540 3012
rect -488 2960 -480 3012
rect -548 2952 -480 2960
rect -402 3012 -334 3022
rect -304 3018 -160 3024
rect -402 2960 -392 3012
rect -340 2960 -334 3012
rect -402 2952 -334 2960
rect 1726 3014 1792 3024
rect 1726 2962 1732 3014
rect 1784 2962 1792 3014
rect 1726 2952 1792 2962
rect -2332 2948 -2188 2952
rect -2332 2946 -2324 2948
rect -2577 2940 -2324 2946
rect -2198 2946 -2188 2948
rect 1306 2946 1316 2948
rect -2198 2940 -578 2946
rect -2577 2906 -2565 2940
rect -590 2906 -578 2940
rect -2577 2900 -2324 2906
rect -2332 2896 -2324 2900
rect -2198 2900 -578 2906
rect -305 2940 1316 2946
rect 1442 2946 1450 2948
rect 1442 2940 1694 2946
rect -305 2906 -293 2940
rect 1682 2906 1694 2940
rect -305 2900 1316 2906
rect -2198 2896 -2188 2900
rect 1306 2896 1316 2900
rect 1442 2900 1694 2906
rect 1442 2896 1450 2900
rect -2332 2890 -2188 2896
rect -3002 2734 -394 2786
rect -342 2734 1734 2786
rect 1786 2734 1792 2786
rect -2334 2654 -2324 2706
rect -2198 2654 1556 2706
rect 1682 2654 1690 2706
rect -2574 2574 -2564 2626
rect -2438 2574 1314 2626
rect 1440 2574 1450 2626
rect -2870 2350 -2780 2402
rect -2004 2398 -1994 2402
rect -2004 2350 -1914 2398
rect -1620 2350 -1610 2402
rect -634 2350 -624 2402
rect -226 2350 -216 2402
rect 760 2350 770 2402
rect 1038 2350 1120 2402
rect 1896 2350 1988 2402
rect -2870 2272 -2824 2350
rect -1960 2330 -1914 2350
rect 1038 2346 1110 2350
rect 1038 2330 1078 2346
rect -1960 2272 -1660 2330
rect -604 2272 -594 2330
rect -2870 2220 -594 2272
rect -2870 2150 -2824 2220
rect -1960 2162 -1660 2220
rect -604 2162 -594 2220
rect -542 2162 -532 2330
rect -318 2162 -308 2330
rect -256 2272 -246 2330
rect 810 2272 1078 2330
rect 1942 2314 1988 2350
rect 1948 2272 1982 2314
rect -256 2220 1988 2272
rect -256 2162 -246 2220
rect 810 2162 1078 2220
rect 1948 2162 1982 2220
rect -1960 2150 -1914 2162
rect -2730 2020 -2056 2134
rect -1472 2020 -798 2140
rect -50 2020 624 2134
rect -3002 1986 2120 2020
rect -3002 1540 -1818 1986
rect -1620 1864 -1610 1916
rect -634 1864 -624 1916
rect -226 1864 -216 1916
rect 760 1864 770 1916
rect -604 1788 -594 1844
rect -1700 1736 -594 1788
rect -604 1676 -594 1736
rect -542 1676 -532 1844
rect -318 1676 -308 1844
rect -256 1788 -246 1844
rect -256 1736 844 1788
rect -256 1676 -246 1736
rect -1610 1540 -634 1648
rect -216 1540 760 1648
rect 936 1540 2120 1986
rect -3002 1534 2120 1540
rect -3002 1500 -2968 1534
rect 2084 1500 2120 1534
rect -3002 1464 2120 1500
rect 936 1462 2120 1464
<< via1 >>
rect -2196 4716 -620 4768
rect -264 4716 1312 4768
rect -1510 4212 -1458 4380
rect 618 4212 670 4380
rect -1407 4144 569 4196
rect -2666 3924 -2614 3976
rect -540 3924 -488 3976
rect -712 3788 -586 3796
rect -712 3754 -590 3788
rect -590 3754 -586 3788
rect -712 3744 -586 3754
rect -296 3788 -170 3796
rect -296 3754 -293 3788
rect -293 3754 -170 3788
rect -296 3744 -170 3754
rect -2564 3660 -2438 3668
rect -2564 3626 -2438 3660
rect -2564 3616 -2438 3626
rect 1556 3660 1682 3668
rect 1556 3626 1682 3660
rect 1556 3616 1682 3626
rect -712 3548 -586 3556
rect -712 3514 -590 3548
rect -590 3514 -586 3548
rect -712 3504 -586 3514
rect -296 3548 -170 3556
rect -296 3514 -293 3548
rect -293 3514 -170 3548
rect -296 3504 -170 3514
rect -2666 3486 -2614 3494
rect -2666 3448 -2658 3486
rect -2658 3448 -2624 3486
rect -2624 3448 -2614 3486
rect -2666 3442 -2614 3448
rect -540 3486 -488 3492
rect -540 3448 -531 3486
rect -531 3448 -497 3486
rect -497 3448 -488 3486
rect -540 3440 -488 3448
rect -392 3486 -340 3492
rect -392 3448 -386 3486
rect -386 3448 -352 3486
rect -352 3448 -340 3486
rect -392 3440 -340 3448
rect 1732 3486 1784 3494
rect 1732 3448 1741 3486
rect 1741 3448 1775 3486
rect 1775 3448 1784 3486
rect 1732 3442 1784 3448
rect -2324 3420 -2198 3428
rect -2324 3386 -2198 3420
rect -2324 3376 -2198 3386
rect 1316 3420 1442 3428
rect 1316 3386 1442 3420
rect 1316 3376 1442 3386
rect -712 3308 -586 3316
rect -712 3274 -590 3308
rect -590 3274 -586 3308
rect -712 3264 -586 3274
rect -296 3308 -170 3316
rect -296 3274 -293 3308
rect -293 3274 -170 3308
rect -296 3264 -170 3274
rect -2564 3180 -2438 3188
rect -2564 3146 -2438 3180
rect -2564 3136 -2438 3146
rect 1556 3180 1682 3188
rect 1556 3146 1682 3180
rect 1556 3136 1682 3146
rect -712 3068 -586 3076
rect -712 3034 -590 3068
rect -590 3034 -586 3068
rect -712 3024 -586 3034
rect -296 3068 -170 3076
rect -296 3034 -293 3068
rect -293 3034 -170 3068
rect -296 3024 -170 3034
rect -2666 3006 -2614 3014
rect -2666 2968 -2658 3006
rect -2658 2968 -2624 3006
rect -2624 2968 -2614 3006
rect -2666 2962 -2614 2968
rect -540 3006 -488 3012
rect -540 2968 -531 3006
rect -531 2968 -497 3006
rect -497 2968 -488 3006
rect -540 2960 -488 2968
rect -392 3006 -340 3012
rect -392 2968 -386 3006
rect -386 2968 -352 3006
rect -352 2968 -340 3006
rect -392 2960 -340 2968
rect 1732 3006 1784 3014
rect 1732 2968 1741 3006
rect 1741 2968 1775 3006
rect 1775 2968 1784 3006
rect 1732 2962 1784 2968
rect -2324 2940 -2198 2948
rect -2324 2906 -2198 2940
rect -2324 2896 -2198 2906
rect 1316 2940 1442 2948
rect 1316 2906 1442 2940
rect 1316 2896 1442 2906
rect -394 2734 -342 2786
rect 1734 2734 1786 2786
rect -2324 2654 -2198 2706
rect 1556 2654 1682 2706
rect -2564 2574 -2438 2626
rect 1314 2574 1440 2626
rect -2780 2350 -2004 2402
rect -1610 2350 -634 2402
rect -216 2350 760 2402
rect 1120 2350 1896 2402
rect -594 2162 -542 2330
rect -308 2162 -256 2330
rect -1610 1864 -634 1916
rect -216 1864 760 1916
rect -594 1676 -542 1844
rect -308 1676 -256 1844
<< metal2 >>
rect -3002 5028 -416 5080
rect -2196 4768 -620 4778
rect -2976 4716 -2196 4768
rect -2976 1916 -2924 4716
rect -2196 4706 -620 4716
rect -1510 4380 -1458 4390
rect -468 4322 -416 5028
rect -264 4768 1312 4778
rect 1312 4716 2120 4768
rect -264 4706 1312 4716
rect 618 4380 670 4390
rect -1458 4270 618 4322
rect -468 4268 -416 4270
rect -1510 4202 -1458 4212
rect -1407 4196 569 4206
rect 618 4202 670 4212
rect -1407 4134 569 4144
rect -722 4037 -160 4134
rect -2674 3924 -2666 3976
rect -2614 3924 -2606 3976
rect -2674 3494 -2606 3924
rect -720 3796 -576 4037
rect -720 3744 -712 3796
rect -586 3744 -576 3796
rect -2674 3442 -2666 3494
rect -2614 3442 -2606 3494
rect -2674 3432 -2606 3442
rect -2572 3668 -2428 3674
rect -2572 3616 -2564 3668
rect -2438 3616 -2428 3668
rect -2674 3022 -2608 3432
rect -2572 3188 -2428 3616
rect -720 3556 -576 3744
rect -720 3504 -712 3556
rect -586 3504 -576 3556
rect -2572 3136 -2564 3188
rect -2438 3136 -2428 3188
rect -2674 3014 -2606 3022
rect -2674 2962 -2666 3014
rect -2614 2962 -2606 3014
rect -2674 2952 -2606 2962
rect -2572 2626 -2428 3136
rect -2332 3428 -2188 3432
rect -2332 3376 -2324 3428
rect -2198 3376 -2188 3428
rect -2332 2948 -2188 3376
rect -720 3316 -576 3504
rect -720 3264 -712 3316
rect -586 3264 -576 3316
rect -720 3076 -576 3264
rect -720 3024 -712 3076
rect -586 3024 -576 3076
rect -720 3022 -576 3024
rect -548 3924 -540 3976
rect -488 3924 -480 3976
rect -548 3492 -480 3924
rect -304 3796 -160 4037
rect -304 3744 -296 3796
rect -170 3744 -160 3796
rect -304 3556 -160 3744
rect -304 3504 -296 3556
rect -170 3504 -160 3556
rect -548 3440 -540 3492
rect -488 3440 -480 3492
rect -548 3012 -480 3440
rect -548 2960 -540 3012
rect -488 2960 -480 3012
rect -548 2952 -480 2960
rect -402 3492 -334 3502
rect -402 3440 -392 3492
rect -340 3440 -334 3492
rect -402 3012 -334 3440
rect -304 3316 -160 3504
rect 1546 3668 1690 3676
rect 1546 3616 1556 3668
rect 1682 3616 1690 3668
rect -304 3264 -296 3316
rect -170 3264 -160 3316
rect -304 3076 -160 3264
rect -304 3024 -296 3076
rect -170 3024 -160 3076
rect -304 3018 -160 3024
rect 1306 3376 1316 3428
rect 1442 3376 1450 3428
rect -402 2960 -392 3012
rect -340 2960 -334 3012
rect -2332 2896 -2324 2948
rect -2198 2896 -2188 2948
rect -2332 2706 -2188 2896
rect -402 2786 -334 2960
rect -402 2734 -394 2786
rect -342 2734 -334 2786
rect 1306 2948 1450 3376
rect 1306 2896 1316 2948
rect 1442 2896 1450 2948
rect -2332 2654 -2324 2706
rect -2198 2654 -2188 2706
rect -2332 2640 -2188 2654
rect -2572 2574 -2564 2626
rect -2438 2574 -2428 2626
rect -2572 2412 -2428 2574
rect -2240 2496 -2188 2640
rect 1306 2626 1450 2896
rect 1306 2574 1314 2626
rect 1440 2574 1450 2626
rect 1546 3188 1690 3616
rect 1546 3136 1556 3188
rect 1682 3136 1690 3188
rect 1546 2706 1690 3136
rect 1726 3494 1792 3504
rect 1726 3442 1732 3494
rect 1784 3442 1792 3494
rect 1726 3014 1792 3442
rect 1726 2962 1732 3014
rect 1784 2962 1792 3014
rect 1726 2786 1792 2962
rect 1726 2734 1734 2786
rect 1786 2734 1792 2786
rect 1546 2654 1556 2706
rect 1682 2654 1690 2706
rect 1306 2564 1440 2574
rect -1610 2496 -1558 2498
rect 1306 2496 1358 2564
rect -2240 2444 -1558 2496
rect -1610 2412 -1558 2444
rect 708 2444 1358 2496
rect 708 2412 760 2444
rect 1546 2412 1690 2654
rect -2780 2402 -2004 2412
rect -2780 2340 -2004 2350
rect -1610 2402 -634 2412
rect -1610 2340 -634 2350
rect -216 2402 760 2412
rect -216 2340 760 2350
rect 1120 2402 1896 2412
rect 1120 2340 1896 2350
rect -594 2330 -542 2340
rect -1610 1916 -634 1926
rect -2976 1864 -1610 1916
rect -1610 1854 -634 1864
rect -594 1844 -542 2162
rect -594 1666 -542 1676
rect -308 2330 -256 2340
rect -308 1844 -256 2162
rect -216 1916 760 1926
rect 2042 1916 2094 4716
rect 760 1864 2094 1916
rect -216 1854 760 1864
rect -308 1666 -256 1676
use sky130_fd_pr__pfet_01v8_lvt_5VNMZ8  sky130_fd_pr__pfet_01v8_lvt_5VNMZ8_0
timestamp 1711036998
transform 0 -1 -1407 1 0 4870
box -296 -1019 296 1019
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_cs_left
timestamp 1711041810
transform 0 -1 -1122 1 0 2246
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_cs_right1
timestamp 1711041810
transform 0 -1 272 1 0 2246
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XMn_diode_left1
timestamp 1711036998
transform 0 -1 -2392 1 0 2246
box -296 -610 296 610
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XMn_diode_right
timestamp 1711036998
transform 0 -1 1510 1 0 2246
box -296 -610 296 610
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_out_left
timestamp 1711041810
transform 0 -1 -1122 1 0 1760
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_out_right
timestamp 1711041810
transform 0 -1 272 1 0 1760
box -296 -734 296 766
use sky130_fd_pr__pfet_01v8_lvt_5VNMZ8  XMp_out
timestamp 1711036998
transform 0 -1 525 1 0 4870
box -296 -1019 296 1019
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_tail
timestamp 1711036998
transform 0 -1 -419 1 0 4296
box -296 -1219 296 1219
<< labels >>
flabel metal1 -2968 5096 2084 5130 0 FreeSans 640 0 0 0 vdd
port 2 nsew default bidirectional
flabel metal2 2068 4716 2120 4768 7 FreeSans 640 0 0 0 vout
port 1 w default output
flabel metal2 -3002 5028 -2950 5080 3 FreeSans 640 0 0 0 vbias_p
port 5 e default input
flabel metal1 -2968 1500 2084 1534 0 FreeSans 640 0 0 0 vss
port 3 nsew default bidirectional
flabel metal1 -3002 3924 -2950 3976 3 FreeSans 640 0 0 0 vinp
port 0 e default input
flabel metal1 -3002 2734 -2950 2786 3 FreeSans 640 0 0 0 vinn
port 4 e default input
flabel metal2 1618 2568 1618 2568 1 FreeSans 320 0 0 0 latch_right
<< end >>
