VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_vaf_555_timer
  CLASS BLOCK ;
  FOREIGN tt_um_vaf_555_timer ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.993000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.993000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 8.700000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 11.400 40.380 18.900 43.250 ;
        RECT 6.080 29.690 18.900 40.380 ;
        RECT 20.375 38.300 45.985 43.690 ;
      LAYER nwell ;
        RECT 6.310 26.470 18.500 29.430 ;
      LAYER pwell ;
        RECT 6.080 18.070 18.900 26.220 ;
      LAYER nwell ;
        RECT 20.375 25.290 45.985 38.300 ;
        RECT 20.370 25.180 45.985 25.290 ;
        RECT 2.725 17.705 9.715 17.710 ;
        RECT 2.725 14.430 19.010 17.705 ;
      LAYER pwell ;
        RECT 2.725 14.425 9.715 14.430 ;
      LAYER nwell ;
        RECT 9.715 14.425 19.010 14.430 ;
      LAYER pwell ;
        RECT 2.725 12.310 19.010 14.425 ;
        RECT 2.725 12.280 4.135 12.310 ;
        RECT 6.320 12.305 19.010 12.310 ;
        RECT 9.715 12.275 19.010 12.305 ;
      LAYER nwell ;
        RECT 20.370 12.170 45.980 25.180 ;
      LAYER pwell ;
        RECT 6.310 7.210 18.410 12.080 ;
        RECT 20.370 6.780 45.980 12.170 ;
      LAYER li1 ;
        RECT 20.545 43.340 45.805 43.510 ;
        RECT 11.580 42.900 18.720 43.070 ;
        RECT 11.580 40.640 11.750 42.900 ;
        RECT 12.630 42.500 17.510 42.900 ;
        RECT 12.550 42.330 17.590 42.500 ;
        RECT 12.210 41.270 12.380 42.270 ;
        RECT 17.760 41.270 17.930 42.270 ;
        RECT 12.550 41.040 17.590 41.210 ;
        RECT 18.550 40.640 18.720 42.900 ;
        RECT 11.580 40.470 18.720 40.640 ;
        RECT 20.545 41.080 26.295 43.340 ;
        RECT 27.255 42.770 32.295 42.940 ;
        RECT 26.915 41.710 27.085 42.710 ;
        RECT 32.465 41.710 32.635 42.710 ;
        RECT 27.255 41.480 32.295 41.650 ;
        RECT 33.095 41.080 33.265 43.340 ;
        RECT 34.225 42.770 39.265 42.940 ;
        RECT 33.885 41.710 34.055 42.710 ;
        RECT 39.435 41.710 39.605 42.710 ;
        RECT 34.225 41.480 39.265 41.650 ;
        RECT 40.065 41.080 45.805 43.340 ;
        RECT 20.545 40.500 45.805 41.080 ;
        RECT 12.180 40.200 17.960 40.470 ;
        RECT 6.260 40.030 18.720 40.200 ;
        RECT 6.260 37.660 6.430 40.030 ;
        RECT 6.910 38.140 9.070 39.550 ;
        RECT 15.910 38.140 18.070 39.550 ;
        RECT 18.550 37.660 18.720 40.030 ;
        RECT 20.555 38.650 20.725 40.500 ;
        RECT 21.405 40.340 25.445 40.500 ;
        RECT 21.485 40.310 25.365 40.340 ;
        RECT 21.065 39.280 21.235 40.280 ;
        RECT 25.615 39.280 25.785 40.280 ;
        RECT 21.405 39.050 25.445 39.220 ;
        RECT 26.125 38.650 26.295 40.500 ;
        RECT 27.255 40.340 32.295 40.500 ;
        RECT 26.915 39.280 27.085 40.280 ;
        RECT 32.465 39.280 32.635 40.280 ;
        RECT 27.255 39.050 32.295 39.220 ;
        RECT 33.095 38.650 33.265 40.500 ;
        RECT 34.225 40.340 39.265 40.500 ;
        RECT 33.885 39.280 34.055 40.280 ;
        RECT 39.435 39.280 39.605 40.280 ;
        RECT 34.225 39.050 39.265 39.220 ;
        RECT 40.065 38.650 40.235 40.500 ;
        RECT 40.915 40.340 44.955 40.500 ;
        RECT 40.995 40.310 44.875 40.340 ;
        RECT 40.575 39.280 40.745 40.280 ;
        RECT 45.125 39.280 45.295 40.280 ;
        RECT 40.915 39.050 44.955 39.220 ;
        RECT 45.635 38.650 45.805 40.500 ;
        RECT 20.555 38.480 45.805 38.650 ;
        RECT 6.260 37.490 18.720 37.660 ;
        RECT 6.260 35.120 6.430 37.490 ;
        RECT 6.910 35.600 9.070 37.010 ;
        RECT 15.910 35.600 18.070 37.010 ;
        RECT 18.550 35.120 18.720 37.490 ;
        RECT 6.260 34.950 18.720 35.120 ;
        RECT 6.260 32.580 6.430 34.950 ;
        RECT 6.910 33.060 9.070 34.470 ;
        RECT 15.910 33.060 18.070 34.470 ;
        RECT 18.550 32.580 18.720 34.950 ;
        RECT 6.260 32.410 18.720 32.580 ;
        RECT 6.260 30.040 6.430 32.410 ;
        RECT 6.910 30.520 9.070 31.930 ;
        RECT 15.910 30.520 18.070 31.930 ;
        RECT 18.550 30.040 18.720 32.410 ;
        RECT 6.260 29.870 18.720 30.040 ;
        RECT 20.545 36.810 45.805 36.980 ;
        RECT 20.545 31.740 21.905 36.810 ;
        RECT 22.480 36.310 32.515 36.480 ;
        RECT 22.095 35.900 22.265 36.250 ;
        RECT 32.730 35.900 32.900 36.250 ;
        RECT 22.480 35.670 32.515 35.840 ;
        RECT 22.480 35.110 32.515 35.280 ;
        RECT 22.095 34.700 22.265 35.050 ;
        RECT 32.730 34.700 32.900 35.050 ;
        RECT 22.480 34.470 32.515 34.640 ;
        RECT 22.480 33.910 32.515 34.080 ;
        RECT 22.095 33.500 22.265 33.850 ;
        RECT 32.730 33.500 32.900 33.850 ;
        RECT 22.480 33.270 32.515 33.440 ;
        RECT 22.480 32.710 32.515 32.880 ;
        RECT 22.095 32.300 22.265 32.650 ;
        RECT 32.730 32.300 32.900 32.650 ;
        RECT 22.480 32.070 32.515 32.240 ;
        RECT 33.095 31.740 33.265 36.810 ;
        RECT 33.840 36.310 43.875 36.480 ;
        RECT 33.455 35.900 33.625 36.250 ;
        RECT 44.090 35.900 44.260 36.250 ;
        RECT 33.840 35.670 43.875 35.840 ;
        RECT 43.115 35.280 43.835 35.370 ;
        RECT 33.840 35.110 43.875 35.280 ;
        RECT 33.455 34.700 33.625 35.050 ;
        RECT 43.115 35.030 43.835 35.110 ;
        RECT 44.090 34.700 44.260 35.050 ;
        RECT 33.840 34.470 43.875 34.640 ;
        RECT 33.840 33.910 43.875 34.080 ;
        RECT 33.455 33.500 33.625 33.850 ;
        RECT 44.090 33.500 44.260 33.850 ;
        RECT 33.840 33.270 43.875 33.440 ;
        RECT 43.115 32.880 43.835 32.970 ;
        RECT 33.840 32.710 43.875 32.880 ;
        RECT 33.455 32.300 33.625 32.650 ;
        RECT 43.115 32.630 43.835 32.710 ;
        RECT 44.090 32.300 44.260 32.650 ;
        RECT 33.840 32.070 43.875 32.240 ;
        RECT 44.450 31.740 45.805 36.810 ;
        RECT 20.545 30.660 45.805 31.740 ;
        RECT 6.490 29.080 18.320 29.250 ;
        RECT 6.490 26.820 6.660 29.080 ;
        RECT 7.385 28.510 17.425 28.680 ;
        RECT 7.000 27.450 7.170 28.450 ;
        RECT 17.640 27.450 17.810 28.450 ;
        RECT 7.385 27.220 17.425 27.390 ;
        RECT 18.150 26.820 18.320 29.080 ;
        RECT 6.490 26.650 18.320 26.820 ;
        RECT 20.545 28.400 27.545 30.660 ;
        RECT 28.270 30.090 38.310 30.260 ;
        RECT 27.885 29.030 28.055 30.030 ;
        RECT 38.525 29.030 38.695 30.030 ;
        RECT 28.270 28.800 38.310 28.970 ;
        RECT 28.350 28.400 38.230 28.800 ;
        RECT 39.025 28.400 45.805 30.660 ;
        RECT 20.545 27.790 45.805 28.400 ;
        RECT 6.260 25.870 18.720 26.040 ;
        RECT 6.260 23.500 6.430 25.870 ;
        RECT 6.910 23.980 9.070 25.390 ;
        RECT 15.910 23.980 18.070 25.390 ;
        RECT 18.550 23.500 18.720 25.870 ;
        RECT 20.545 25.530 23.615 27.790 ;
        RECT 24.330 27.220 32.370 27.390 ;
        RECT 23.945 26.160 24.115 27.160 ;
        RECT 32.585 26.160 32.755 27.160 ;
        RECT 24.330 25.930 32.370 26.100 ;
        RECT 33.095 25.530 33.265 27.790 ;
        RECT 39.025 27.780 45.805 27.790 ;
        RECT 33.990 27.220 42.030 27.390 ;
        RECT 33.605 26.160 33.775 27.160 ;
        RECT 42.245 26.160 42.415 27.160 ;
        RECT 33.990 25.930 42.030 26.100 ;
        RECT 42.755 25.530 45.805 27.780 ;
        RECT 20.545 25.360 45.805 25.530 ;
        RECT 6.260 23.330 18.720 23.500 ;
        RECT 6.260 20.960 6.430 23.330 ;
        RECT 6.910 21.440 9.070 22.850 ;
        RECT 15.910 21.440 18.070 22.850 ;
        RECT 18.550 20.960 18.720 23.330 ;
        RECT 6.260 20.790 18.720 20.960 ;
        RECT 6.260 18.420 6.430 20.790 ;
        RECT 6.910 18.900 9.070 20.310 ;
        RECT 15.910 18.900 18.070 20.310 ;
        RECT 18.550 18.420 18.720 20.790 ;
        RECT 6.260 18.250 18.720 18.420 ;
        RECT 20.540 24.940 45.800 25.110 ;
        RECT 20.540 22.680 23.610 24.940 ;
        RECT 24.325 24.370 32.365 24.540 ;
        RECT 23.940 23.310 24.110 24.310 ;
        RECT 32.580 23.310 32.750 24.310 ;
        RECT 24.325 23.080 32.365 23.250 ;
        RECT 33.090 22.680 33.260 24.940 ;
        RECT 33.985 24.370 42.025 24.540 ;
        RECT 33.600 23.310 33.770 24.310 ;
        RECT 42.240 23.310 42.410 24.310 ;
        RECT 33.985 23.080 42.025 23.250 ;
        RECT 42.750 22.690 45.800 24.940 ;
        RECT 39.020 22.680 45.800 22.690 ;
        RECT 20.540 22.070 45.800 22.680 ;
        RECT 20.540 19.810 27.540 22.070 ;
        RECT 28.345 21.670 38.225 22.070 ;
        RECT 28.265 21.500 38.305 21.670 ;
        RECT 27.880 20.440 28.050 21.440 ;
        RECT 38.520 20.440 38.690 21.440 ;
        RECT 28.265 20.210 38.305 20.380 ;
        RECT 39.020 19.810 45.800 22.070 ;
        RECT 20.540 18.730 45.800 19.810 ;
        RECT 2.725 17.360 4.135 17.530 ;
        RECT 4.365 17.360 5.715 17.530 ;
        RECT 6.220 17.360 7.570 17.530 ;
        RECT 8.100 17.360 9.450 17.530 ;
        RECT 3.125 16.070 3.295 17.110 ;
        RECT 3.565 16.070 3.735 17.110 ;
        RECT 3.265 15.685 3.595 15.855 ;
        RECT 4.495 14.950 4.665 16.990 ;
        RECT 4.935 14.950 5.105 17.360 ;
        RECT 9.715 17.355 19.010 17.525 ;
        RECT 5.375 14.950 5.545 16.990 ;
        RECT 6.355 14.950 6.525 16.990 ;
        RECT 6.795 14.950 6.965 16.990 ;
        RECT 7.235 14.950 7.405 16.990 ;
        RECT 8.235 14.950 8.405 16.990 ;
        RECT 8.675 14.950 8.845 16.990 ;
        RECT 9.115 14.950 9.285 16.990 ;
        RECT 10.115 16.065 10.285 17.105 ;
        RECT 10.555 16.065 10.725 17.105 ;
        RECT 11.425 16.065 11.595 17.105 ;
        RECT 11.865 16.065 12.035 17.105 ;
        RECT 12.740 16.065 12.910 17.105 ;
        RECT 13.180 16.065 13.350 17.105 ;
        RECT 14.055 16.065 14.225 17.105 ;
        RECT 14.495 16.065 14.665 17.105 ;
        RECT 15.370 16.065 15.540 17.105 ;
        RECT 15.810 16.065 15.980 17.105 ;
        RECT 16.685 16.065 16.855 17.105 ;
        RECT 17.125 16.065 17.295 17.105 ;
        RECT 18.000 16.065 18.170 17.105 ;
        RECT 18.440 16.065 18.610 17.105 ;
        RECT 10.255 15.680 10.585 15.850 ;
        RECT 11.565 15.680 11.895 15.850 ;
        RECT 12.880 15.680 13.210 15.850 ;
        RECT 14.195 15.680 14.525 15.850 ;
        RECT 15.510 15.680 15.840 15.850 ;
        RECT 16.825 15.680 17.155 15.850 ;
        RECT 18.140 15.680 18.470 15.850 ;
        RECT 4.535 14.375 4.865 14.705 ;
        RECT 6.480 14.565 6.810 14.735 ;
        RECT 8.360 14.565 8.690 14.735 ;
        RECT 6.580 14.470 6.750 14.565 ;
        RECT 8.460 14.470 8.630 14.565 ;
        RECT 3.265 14.015 3.595 14.185 ;
        RECT 5.085 14.035 5.415 14.205 ;
        RECT 6.940 14.035 7.270 14.205 ;
        RECT 8.820 14.035 9.150 14.205 ;
        RECT 5.185 13.940 5.355 14.035 ;
        RECT 7.040 13.940 7.210 14.035 ;
        RECT 8.920 13.940 9.090 14.035 ;
        RECT 10.255 14.010 10.585 14.180 ;
        RECT 11.565 14.010 11.895 14.180 ;
        RECT 12.880 14.010 13.210 14.180 ;
        RECT 14.195 14.010 14.525 14.180 ;
        RECT 15.510 14.010 15.840 14.180 ;
        RECT 16.825 14.010 17.155 14.180 ;
        RECT 18.140 14.010 18.470 14.180 ;
        RECT 3.125 12.730 3.295 13.770 ;
        RECT 3.565 13.690 3.735 13.770 ;
        RECT 3.555 12.725 3.745 13.690 ;
        RECT 4.495 12.730 4.665 13.770 ;
        RECT 4.935 12.720 5.105 13.770 ;
        RECT 5.375 13.690 5.545 13.770 ;
        RECT 5.365 12.725 5.555 13.690 ;
        RECT 6.350 12.730 6.520 13.770 ;
        RECT 6.790 12.480 6.960 13.770 ;
        RECT 7.230 13.690 7.400 13.770 ;
        RECT 7.220 12.725 7.410 13.690 ;
        RECT 8.230 12.730 8.400 13.770 ;
        RECT 8.670 12.480 8.840 13.770 ;
        RECT 9.110 13.690 9.280 13.770 ;
        RECT 9.100 12.725 9.290 13.690 ;
        RECT 10.115 12.725 10.285 13.765 ;
        RECT 10.555 13.685 10.725 13.765 ;
        RECT 10.545 12.720 10.735 13.685 ;
        RECT 11.425 12.725 11.595 13.765 ;
        RECT 11.865 13.685 12.035 13.765 ;
        RECT 11.855 12.720 12.045 13.685 ;
        RECT 12.740 12.725 12.910 13.765 ;
        RECT 13.180 13.685 13.350 13.765 ;
        RECT 13.170 12.720 13.360 13.685 ;
        RECT 14.055 12.725 14.225 13.765 ;
        RECT 14.495 13.685 14.665 13.765 ;
        RECT 14.485 12.720 14.675 13.685 ;
        RECT 15.370 12.725 15.540 13.765 ;
        RECT 15.810 13.685 15.980 13.765 ;
        RECT 15.800 12.720 15.990 13.685 ;
        RECT 16.685 12.725 16.855 13.765 ;
        RECT 17.125 13.685 17.295 13.765 ;
        RECT 17.115 12.720 17.305 13.685 ;
        RECT 18.000 12.725 18.170 13.765 ;
        RECT 18.440 13.685 18.610 13.765 ;
        RECT 18.430 12.720 18.620 13.685 ;
        RECT 20.540 13.660 21.900 18.730 ;
        RECT 22.475 18.230 32.510 18.400 ;
        RECT 22.090 17.820 22.260 18.170 ;
        RECT 32.725 17.820 32.895 18.170 ;
        RECT 22.475 17.590 32.510 17.760 ;
        RECT 22.475 17.030 32.510 17.200 ;
        RECT 22.090 16.620 22.260 16.970 ;
        RECT 32.725 16.620 32.895 16.970 ;
        RECT 22.475 16.390 32.510 16.560 ;
        RECT 22.475 15.830 32.510 16.000 ;
        RECT 22.090 15.420 22.260 15.770 ;
        RECT 32.725 15.420 32.895 15.770 ;
        RECT 22.475 15.190 32.510 15.360 ;
        RECT 22.475 14.630 32.510 14.800 ;
        RECT 22.090 14.220 22.260 14.570 ;
        RECT 32.725 14.220 32.895 14.570 ;
        RECT 22.475 13.990 32.510 14.160 ;
        RECT 33.090 13.660 33.260 18.730 ;
        RECT 33.835 18.230 43.870 18.400 ;
        RECT 33.450 17.820 33.620 18.170 ;
        RECT 43.110 17.760 43.830 17.840 ;
        RECT 44.085 17.820 44.255 18.170 ;
        RECT 33.835 17.590 43.870 17.760 ;
        RECT 43.110 17.500 43.830 17.590 ;
        RECT 33.835 17.030 43.870 17.200 ;
        RECT 33.450 16.620 33.620 16.970 ;
        RECT 44.085 16.620 44.255 16.970 ;
        RECT 33.835 16.390 43.870 16.560 ;
        RECT 33.835 15.830 43.870 16.000 ;
        RECT 33.450 15.420 33.620 15.770 ;
        RECT 43.110 15.360 43.830 15.440 ;
        RECT 44.085 15.420 44.255 15.770 ;
        RECT 33.835 15.190 43.870 15.360 ;
        RECT 43.110 15.100 43.830 15.190 ;
        RECT 33.835 14.630 43.870 14.800 ;
        RECT 33.450 14.220 33.620 14.570 ;
        RECT 44.085 14.220 44.255 14.570 ;
        RECT 33.835 13.990 43.870 14.160 ;
        RECT 44.445 13.660 45.800 18.730 ;
        RECT 20.540 13.490 45.800 13.660 ;
        RECT 2.915 12.475 9.495 12.480 ;
        RECT 2.915 12.310 18.780 12.475 ;
        RECT 6.315 12.305 18.780 12.310 ;
        RECT 6.315 11.730 18.700 12.305 ;
        RECT 20.550 11.820 45.800 11.990 ;
        RECT 6.490 11.420 6.660 11.730 ;
        RECT 6.400 7.870 6.660 11.420 ;
        RECT 7.340 11.160 17.380 11.330 ;
        RECT 7.000 10.750 7.170 11.100 ;
        RECT 17.550 10.750 17.720 11.100 ;
        RECT 7.340 10.520 17.380 10.690 ;
        RECT 7.000 10.110 7.170 10.460 ;
        RECT 17.550 10.110 17.720 10.460 ;
        RECT 7.340 9.880 17.380 10.050 ;
        RECT 7.000 9.470 7.170 9.820 ;
        RECT 17.550 9.470 17.720 9.820 ;
        RECT 7.340 9.240 17.380 9.410 ;
        RECT 7.000 8.830 7.170 9.180 ;
        RECT 17.550 8.830 17.720 9.180 ;
        RECT 7.340 8.600 17.380 8.770 ;
        RECT 7.000 8.190 7.170 8.540 ;
        RECT 17.550 8.190 17.720 8.540 ;
        RECT 7.340 7.960 17.380 8.130 ;
        RECT 6.490 7.560 6.660 7.870 ;
        RECT 18.060 7.560 18.230 11.730 ;
        RECT 20.550 9.970 20.720 11.820 ;
        RECT 21.400 11.250 25.440 11.420 ;
        RECT 21.060 10.190 21.230 11.190 ;
        RECT 25.610 10.190 25.780 11.190 ;
        RECT 21.480 10.130 25.360 10.160 ;
        RECT 21.400 9.970 25.440 10.130 ;
        RECT 26.120 9.970 26.290 11.820 ;
        RECT 27.250 11.250 32.290 11.420 ;
        RECT 26.910 10.190 27.080 11.190 ;
        RECT 32.460 10.190 32.630 11.190 ;
        RECT 27.250 9.970 32.290 10.130 ;
        RECT 33.090 9.970 33.260 11.820 ;
        RECT 34.220 11.250 39.260 11.420 ;
        RECT 33.880 10.190 34.050 11.190 ;
        RECT 39.430 10.190 39.600 11.190 ;
        RECT 34.220 9.970 39.260 10.130 ;
        RECT 40.060 9.970 40.230 11.820 ;
        RECT 40.910 11.250 44.950 11.420 ;
        RECT 40.570 10.190 40.740 11.190 ;
        RECT 45.120 10.190 45.290 11.190 ;
        RECT 40.990 10.130 44.870 10.160 ;
        RECT 40.910 9.970 44.950 10.130 ;
        RECT 45.630 9.970 45.800 11.820 ;
        RECT 6.490 7.390 18.230 7.560 ;
        RECT 20.540 9.390 45.800 9.970 ;
        RECT 20.540 7.130 26.290 9.390 ;
        RECT 27.250 8.820 32.290 8.990 ;
        RECT 26.910 7.760 27.080 8.760 ;
        RECT 32.460 7.760 32.630 8.760 ;
        RECT 27.250 7.530 32.290 7.700 ;
        RECT 33.090 7.130 33.260 9.390 ;
        RECT 34.220 8.820 39.260 8.990 ;
        RECT 33.880 7.760 34.050 8.760 ;
        RECT 39.430 7.760 39.600 8.760 ;
        RECT 34.220 7.530 39.260 7.700 ;
        RECT 40.060 7.130 45.800 9.390 ;
        RECT 20.540 6.960 45.800 7.130 ;
      LAYER mcon ;
        RECT 20.545 43.340 45.805 43.510 ;
        RECT 12.630 42.330 17.510 42.500 ;
        RECT 12.210 41.350 12.380 42.190 ;
        RECT 17.760 41.350 17.930 42.190 ;
        RECT 12.630 41.040 17.510 41.210 ;
        RECT 27.335 42.770 32.215 42.940 ;
        RECT 26.915 41.790 27.085 42.630 ;
        RECT 32.465 41.790 32.635 42.630 ;
        RECT 27.335 41.480 32.215 41.650 ;
        RECT 34.305 42.770 39.185 42.940 ;
        RECT 33.885 41.790 34.055 42.630 ;
        RECT 39.435 41.790 39.605 42.630 ;
        RECT 34.305 41.480 39.185 41.650 ;
        RECT 7.000 38.220 8.985 39.470 ;
        RECT 15.995 38.220 17.980 39.470 ;
        RECT 21.485 40.340 25.365 40.510 ;
        RECT 21.065 39.360 21.235 40.200 ;
        RECT 25.615 39.360 25.785 40.200 ;
        RECT 21.485 39.050 25.365 39.220 ;
        RECT 27.335 40.340 32.215 40.510 ;
        RECT 26.915 39.360 27.085 40.200 ;
        RECT 32.465 39.360 32.635 40.200 ;
        RECT 27.335 39.050 32.215 39.220 ;
        RECT 34.305 40.340 39.185 40.510 ;
        RECT 33.885 39.360 34.055 40.200 ;
        RECT 39.435 39.360 39.605 40.200 ;
        RECT 34.305 39.050 39.185 39.220 ;
        RECT 40.995 40.340 44.875 40.510 ;
        RECT 40.575 39.360 40.745 40.200 ;
        RECT 45.125 39.360 45.295 40.200 ;
        RECT 40.995 39.050 44.875 39.220 ;
        RECT 7.000 35.680 8.985 36.930 ;
        RECT 15.995 35.680 17.980 36.930 ;
        RECT 7.000 33.140 8.985 34.390 ;
        RECT 15.995 33.140 17.980 34.390 ;
        RECT 7.000 30.600 8.985 31.850 ;
        RECT 15.995 30.600 17.980 31.850 ;
        RECT 22.560 36.310 32.435 36.480 ;
        RECT 22.095 35.980 22.265 36.170 ;
        RECT 32.730 35.980 32.900 36.170 ;
        RECT 22.560 35.670 32.435 35.840 ;
        RECT 22.560 35.110 32.435 35.280 ;
        RECT 22.095 34.780 22.265 34.970 ;
        RECT 32.730 34.780 32.900 34.970 ;
        RECT 22.560 34.470 32.435 34.640 ;
        RECT 22.560 33.910 32.435 34.080 ;
        RECT 22.095 33.580 22.265 33.770 ;
        RECT 32.730 33.580 32.900 33.770 ;
        RECT 22.560 33.270 32.435 33.440 ;
        RECT 22.560 32.710 32.435 32.880 ;
        RECT 22.095 32.380 22.265 32.570 ;
        RECT 32.730 32.380 32.900 32.570 ;
        RECT 22.560 32.070 32.435 32.240 ;
        RECT 33.920 36.310 43.795 36.480 ;
        RECT 33.455 35.980 33.625 36.170 ;
        RECT 44.090 35.980 44.260 36.170 ;
        RECT 33.920 35.670 43.795 35.840 ;
        RECT 33.920 35.110 43.815 35.280 ;
        RECT 33.455 34.780 33.625 34.970 ;
        RECT 44.090 34.780 44.260 34.970 ;
        RECT 33.920 34.470 43.795 34.640 ;
        RECT 33.920 33.910 43.795 34.080 ;
        RECT 33.455 33.580 33.625 33.770 ;
        RECT 44.090 33.580 44.260 33.770 ;
        RECT 33.920 33.270 43.795 33.440 ;
        RECT 33.920 32.710 43.815 32.880 ;
        RECT 33.455 32.380 33.625 32.570 ;
        RECT 44.090 32.380 44.260 32.570 ;
        RECT 33.920 32.070 43.795 32.240 ;
        RECT 7.465 28.510 17.345 28.680 ;
        RECT 7.000 27.530 7.170 28.370 ;
        RECT 17.640 27.530 17.810 28.370 ;
        RECT 7.465 27.220 17.345 27.390 ;
        RECT 6.970 26.650 17.840 26.820 ;
        RECT 28.350 30.090 38.230 30.260 ;
        RECT 27.885 29.110 28.055 29.950 ;
        RECT 38.525 29.110 38.695 29.950 ;
        RECT 28.350 28.800 38.230 28.970 ;
        RECT 7.000 24.060 8.985 25.310 ;
        RECT 15.995 24.060 17.980 25.310 ;
        RECT 24.410 27.220 32.290 27.390 ;
        RECT 23.945 26.240 24.115 27.080 ;
        RECT 32.585 26.240 32.755 27.080 ;
        RECT 24.410 25.930 32.290 26.100 ;
        RECT 34.070 27.220 41.950 27.390 ;
        RECT 33.605 26.240 33.775 27.080 ;
        RECT 42.245 26.240 42.415 27.080 ;
        RECT 34.070 25.930 41.950 26.100 ;
        RECT 20.545 25.360 45.805 25.530 ;
        RECT 7.000 21.520 8.985 22.770 ;
        RECT 15.995 21.520 17.980 22.770 ;
        RECT 7.000 18.980 8.985 20.230 ;
        RECT 15.995 18.980 17.980 20.230 ;
        RECT 20.540 24.940 45.800 25.110 ;
        RECT 24.405 24.370 32.285 24.540 ;
        RECT 23.940 23.390 24.110 24.230 ;
        RECT 32.580 23.390 32.750 24.230 ;
        RECT 24.405 23.080 32.285 23.250 ;
        RECT 34.065 24.370 41.945 24.540 ;
        RECT 33.600 23.390 33.770 24.230 ;
        RECT 42.240 23.390 42.410 24.230 ;
        RECT 34.065 23.080 41.945 23.250 ;
        RECT 28.345 21.500 38.225 21.670 ;
        RECT 27.880 20.520 28.050 21.360 ;
        RECT 38.520 20.520 38.690 21.360 ;
        RECT 28.345 20.210 38.225 20.380 ;
        RECT 3.035 17.360 3.825 17.530 ;
        RECT 4.445 17.360 5.635 17.530 ;
        RECT 6.300 17.360 7.490 17.530 ;
        RECT 8.180 17.360 9.370 17.530 ;
        RECT 3.125 16.150 3.295 17.030 ;
        RECT 3.565 16.150 3.735 17.030 ;
        RECT 3.345 15.685 3.515 15.855 ;
        RECT 4.495 15.030 4.665 16.910 ;
        RECT 10.025 17.355 10.815 17.525 ;
        RECT 11.335 17.355 12.125 17.525 ;
        RECT 12.650 17.355 13.440 17.525 ;
        RECT 13.965 17.355 14.755 17.525 ;
        RECT 15.280 17.355 16.070 17.525 ;
        RECT 16.595 17.355 17.385 17.525 ;
        RECT 17.910 17.355 18.700 17.525 ;
        RECT 5.375 15.030 5.545 16.910 ;
        RECT 6.355 15.030 6.525 16.910 ;
        RECT 7.235 15.030 7.405 16.910 ;
        RECT 8.235 15.030 8.405 16.910 ;
        RECT 9.115 15.030 9.285 16.910 ;
        RECT 10.115 16.145 10.285 17.025 ;
        RECT 10.555 16.145 10.725 17.025 ;
        RECT 11.425 16.145 11.595 17.025 ;
        RECT 11.865 16.145 12.035 17.025 ;
        RECT 12.740 16.145 12.910 17.025 ;
        RECT 13.180 16.145 13.350 17.025 ;
        RECT 14.055 16.145 14.225 17.025 ;
        RECT 14.495 16.145 14.665 17.025 ;
        RECT 15.370 16.145 15.540 17.025 ;
        RECT 15.810 16.145 15.980 17.025 ;
        RECT 16.685 16.145 16.855 17.025 ;
        RECT 17.125 16.145 17.295 17.025 ;
        RECT 18.000 16.145 18.170 17.025 ;
        RECT 18.440 16.145 18.610 17.025 ;
        RECT 10.335 15.680 10.505 15.850 ;
        RECT 11.645 15.680 11.815 15.850 ;
        RECT 12.960 15.680 13.130 15.850 ;
        RECT 14.275 15.680 14.445 15.850 ;
        RECT 15.590 15.680 15.760 15.850 ;
        RECT 16.905 15.680 17.075 15.850 ;
        RECT 18.220 15.680 18.390 15.850 ;
        RECT 4.615 14.455 4.785 14.625 ;
        RECT 6.560 14.565 6.730 14.735 ;
        RECT 8.440 14.565 8.610 14.735 ;
        RECT 3.345 14.015 3.515 14.185 ;
        RECT 5.165 14.035 5.335 14.205 ;
        RECT 7.020 14.035 7.190 14.205 ;
        RECT 8.900 14.035 9.070 14.205 ;
        RECT 10.335 14.010 10.505 14.180 ;
        RECT 11.645 14.010 11.815 14.180 ;
        RECT 12.960 14.010 13.130 14.180 ;
        RECT 14.275 14.010 14.445 14.180 ;
        RECT 15.590 14.010 15.760 14.180 ;
        RECT 16.905 14.010 17.075 14.180 ;
        RECT 18.220 14.010 18.390 14.180 ;
        RECT 3.125 12.810 3.295 13.690 ;
        RECT 3.565 12.805 3.735 13.690 ;
        RECT 4.495 12.810 4.665 13.690 ;
        RECT 5.375 12.805 5.545 13.690 ;
        RECT 6.350 12.810 6.520 13.690 ;
        RECT 7.230 12.805 7.400 13.690 ;
        RECT 8.230 12.810 8.400 13.690 ;
        RECT 9.110 12.805 9.280 13.690 ;
        RECT 10.115 12.805 10.285 13.685 ;
        RECT 10.555 12.800 10.725 13.685 ;
        RECT 11.425 12.805 11.595 13.685 ;
        RECT 11.865 12.800 12.035 13.685 ;
        RECT 12.740 12.805 12.910 13.685 ;
        RECT 13.180 12.800 13.350 13.685 ;
        RECT 14.055 12.805 14.225 13.685 ;
        RECT 14.495 12.800 14.665 13.685 ;
        RECT 15.370 12.805 15.540 13.685 ;
        RECT 15.810 12.800 15.980 13.685 ;
        RECT 16.685 12.805 16.855 13.685 ;
        RECT 17.125 12.800 17.295 13.685 ;
        RECT 18.000 12.805 18.170 13.685 ;
        RECT 18.440 12.800 18.610 13.685 ;
        RECT 22.555 18.230 32.430 18.400 ;
        RECT 22.090 17.900 22.260 18.090 ;
        RECT 32.725 17.900 32.895 18.090 ;
        RECT 22.555 17.590 32.430 17.760 ;
        RECT 22.555 17.030 32.430 17.200 ;
        RECT 22.090 16.700 22.260 16.890 ;
        RECT 32.725 16.700 32.895 16.890 ;
        RECT 22.555 16.390 32.430 16.560 ;
        RECT 22.555 15.830 32.430 16.000 ;
        RECT 22.090 15.500 22.260 15.690 ;
        RECT 32.725 15.500 32.895 15.690 ;
        RECT 22.555 15.190 32.430 15.360 ;
        RECT 22.555 14.630 32.430 14.800 ;
        RECT 22.090 14.300 22.260 14.490 ;
        RECT 32.725 14.300 32.895 14.490 ;
        RECT 22.555 13.990 32.430 14.160 ;
        RECT 33.915 18.230 43.790 18.400 ;
        RECT 33.450 17.900 33.620 18.090 ;
        RECT 44.085 17.900 44.255 18.090 ;
        RECT 33.915 17.590 43.810 17.760 ;
        RECT 33.915 17.030 43.790 17.200 ;
        RECT 33.450 16.700 33.620 16.890 ;
        RECT 44.085 16.700 44.255 16.890 ;
        RECT 33.915 16.390 43.790 16.560 ;
        RECT 33.915 15.830 43.790 16.000 ;
        RECT 33.450 15.500 33.620 15.690 ;
        RECT 44.085 15.500 44.255 15.690 ;
        RECT 33.915 15.190 43.810 15.360 ;
        RECT 33.915 14.630 43.790 14.800 ;
        RECT 33.450 14.300 33.620 14.490 ;
        RECT 44.085 14.300 44.255 14.490 ;
        RECT 33.915 13.990 43.790 14.160 ;
        RECT 3.035 12.310 3.825 12.480 ;
        RECT 4.405 12.310 5.635 12.480 ;
        RECT 6.260 12.310 7.490 12.480 ;
        RECT 8.140 12.310 9.370 12.480 ;
        RECT 10.025 12.305 10.815 12.475 ;
        RECT 11.335 12.305 12.125 12.475 ;
        RECT 12.650 12.305 13.440 12.475 ;
        RECT 13.965 12.305 14.755 12.475 ;
        RECT 15.280 12.305 16.070 12.475 ;
        RECT 16.595 12.305 17.385 12.475 ;
        RECT 17.910 12.305 18.700 12.475 ;
        RECT 6.970 11.730 17.750 11.900 ;
        RECT 6.400 7.870 6.660 11.420 ;
        RECT 7.420 11.160 17.300 11.330 ;
        RECT 7.000 10.830 7.170 11.020 ;
        RECT 17.550 10.830 17.720 11.020 ;
        RECT 7.420 10.520 17.300 10.690 ;
        RECT 7.000 10.190 7.170 10.380 ;
        RECT 17.550 10.190 17.720 10.380 ;
        RECT 7.420 9.880 17.300 10.050 ;
        RECT 7.000 9.550 7.170 9.740 ;
        RECT 17.550 9.550 17.720 9.740 ;
        RECT 7.420 9.240 17.300 9.410 ;
        RECT 7.000 8.910 7.170 9.100 ;
        RECT 17.550 8.910 17.720 9.100 ;
        RECT 7.420 8.600 17.300 8.770 ;
        RECT 7.000 8.270 7.170 8.460 ;
        RECT 17.550 8.270 17.720 8.460 ;
        RECT 7.420 7.960 17.300 8.130 ;
        RECT 21.480 11.250 25.360 11.420 ;
        RECT 21.060 10.270 21.230 11.110 ;
        RECT 25.610 10.270 25.780 11.110 ;
        RECT 21.480 9.960 25.360 10.130 ;
        RECT 27.330 11.250 32.210 11.420 ;
        RECT 26.910 10.270 27.080 11.110 ;
        RECT 32.460 10.270 32.630 11.110 ;
        RECT 27.330 9.960 32.210 10.130 ;
        RECT 34.300 11.250 39.180 11.420 ;
        RECT 33.880 10.270 34.050 11.110 ;
        RECT 39.430 10.270 39.600 11.110 ;
        RECT 34.300 9.960 39.180 10.130 ;
        RECT 40.990 11.250 44.870 11.420 ;
        RECT 40.570 10.270 40.740 11.110 ;
        RECT 45.120 10.270 45.290 11.110 ;
        RECT 40.990 9.960 44.870 10.130 ;
        RECT 27.330 8.820 32.210 8.990 ;
        RECT 26.910 7.840 27.080 8.680 ;
        RECT 32.460 7.840 32.630 8.680 ;
        RECT 27.330 7.530 32.210 7.700 ;
        RECT 34.300 8.820 39.180 8.990 ;
        RECT 33.880 7.840 34.050 8.680 ;
        RECT 39.430 7.840 39.600 8.680 ;
        RECT 34.300 7.530 39.180 7.700 ;
        RECT 20.540 6.960 45.800 7.130 ;
      LAYER met1 ;
        RECT 5.180 50.840 5.550 52.070 ;
        RECT 7.060 50.940 7.430 52.170 ;
        RECT 18.470 46.690 20.580 46.950 ;
        RECT 12.580 42.530 17.560 42.610 ;
        RECT 12.570 42.300 17.570 42.530 ;
        RECT 12.180 41.290 12.410 42.250 ;
        RECT 17.730 41.350 17.960 42.250 ;
        RECT 17.730 41.260 18.070 41.350 ;
        RECT 15.910 41.240 18.070 41.260 ;
        RECT 12.570 41.010 18.070 41.240 ;
        RECT 6.910 35.600 9.070 39.550 ;
        RECT 15.910 38.140 18.070 41.010 ;
        RECT 6.910 30.520 9.070 34.470 ;
        RECT 15.910 33.060 18.070 37.010 ;
        RECT 15.910 28.710 18.070 31.930 ;
        RECT 18.520 31.390 18.780 46.690 ;
        RECT 19.570 45.740 24.160 46.000 ;
        RECT 19.570 41.870 19.830 45.740 ;
        RECT 22.100 45.630 22.360 45.740 ;
        RECT 40.065 43.690 45.985 43.700 ;
        RECT 20.375 43.310 45.985 43.690 ;
        RECT 19.520 41.610 19.880 41.870 ;
        RECT 20.375 41.080 26.295 43.310 ;
        RECT 27.335 42.970 32.215 43.310 ;
        RECT 34.305 42.970 39.185 43.310 ;
        RECT 27.275 42.740 32.275 42.970 ;
        RECT 34.245 42.740 39.245 42.970 ;
        RECT 26.885 42.330 27.115 42.690 ;
        RECT 32.435 42.630 32.665 42.690 ;
        RECT 33.855 42.630 34.085 42.690 ;
        RECT 32.365 42.330 32.725 42.630 ;
        RECT 26.885 42.070 32.725 42.330 ;
        RECT 26.885 41.730 27.115 42.070 ;
        RECT 32.365 41.790 32.725 42.070 ;
        RECT 33.795 42.330 34.155 42.630 ;
        RECT 39.405 42.330 39.635 42.690 ;
        RECT 33.795 42.070 39.635 42.330 ;
        RECT 33.795 41.790 34.155 42.070 ;
        RECT 32.435 41.730 32.665 41.790 ;
        RECT 33.855 41.730 34.085 41.790 ;
        RECT 39.405 41.730 39.635 42.070 ;
        RECT 27.285 41.680 32.265 41.690 ;
        RECT 34.255 41.680 39.235 41.690 ;
        RECT 27.275 41.450 32.275 41.680 ;
        RECT 34.245 41.450 39.245 41.680 ;
        RECT 27.285 41.430 32.265 41.450 ;
        RECT 34.255 41.430 39.235 41.450 ;
        RECT 40.065 41.080 45.985 43.310 ;
        RECT 20.375 40.910 45.985 41.080 ;
        RECT 21.735 40.540 25.105 40.910 ;
        RECT 28.025 40.540 31.395 40.910 ;
        RECT 35.135 40.540 38.505 40.910 ;
        RECT 21.425 40.310 25.425 40.540 ;
        RECT 27.275 40.310 32.275 40.540 ;
        RECT 34.245 40.310 39.245 40.540 ;
        RECT 40.935 40.310 44.935 40.540 ;
        RECT 21.035 39.910 21.265 40.260 ;
        RECT 25.585 40.200 25.815 40.260 ;
        RECT 26.885 40.200 27.115 40.260 ;
        RECT 32.435 40.200 32.665 40.260 ;
        RECT 33.855 40.200 34.085 40.260 ;
        RECT 39.405 40.200 39.635 40.260 ;
        RECT 40.545 40.200 40.775 40.260 ;
        RECT 25.585 39.910 27.115 40.200 ;
        RECT 32.365 39.910 32.725 40.200 ;
        RECT 21.035 39.650 32.725 39.910 ;
        RECT 21.035 39.260 21.265 39.650 ;
        RECT 25.585 39.360 27.115 39.650 ;
        RECT 32.365 39.360 32.725 39.650 ;
        RECT 33.795 39.910 34.155 40.200 ;
        RECT 39.405 39.910 40.775 40.200 ;
        RECT 45.095 39.910 45.325 40.260 ;
        RECT 33.795 39.650 45.325 39.910 ;
        RECT 33.795 39.360 34.155 39.650 ;
        RECT 39.405 39.360 40.775 39.650 ;
        RECT 25.585 39.260 25.815 39.360 ;
        RECT 26.885 39.300 27.115 39.360 ;
        RECT 32.435 39.300 32.665 39.360 ;
        RECT 33.855 39.300 34.085 39.360 ;
        RECT 39.405 39.300 39.635 39.360 ;
        RECT 40.545 39.300 40.775 39.360 ;
        RECT 40.575 39.280 40.775 39.300 ;
        RECT 40.575 39.260 40.935 39.280 ;
        RECT 45.095 39.260 45.325 39.650 ;
        RECT 21.035 39.020 25.815 39.260 ;
        RECT 27.285 39.250 32.265 39.260 ;
        RECT 34.255 39.250 39.235 39.260 ;
        RECT 27.275 39.020 32.275 39.250 ;
        RECT 34.245 39.020 39.245 39.250 ;
        RECT 21.035 39.000 25.415 39.020 ;
        RECT 27.285 39.000 32.265 39.020 ;
        RECT 34.255 39.000 39.235 39.020 ;
        RECT 40.575 39.000 45.325 39.260 ;
        RECT 22.515 37.880 42.635 38.140 ;
        RECT 23.715 37.480 43.835 37.740 ;
        RECT 19.150 37.345 19.530 37.390 ;
        RECT 19.150 37.340 20.410 37.345 ;
        RECT 19.150 37.085 44.345 37.340 ;
        RECT 19.150 37.040 19.530 37.085 ;
        RECT 20.375 37.080 44.345 37.085 ;
        RECT 21.695 34.970 21.885 37.080 ;
        RECT 23.725 36.510 24.445 36.560 ;
        RECT 41.915 36.510 42.635 36.530 ;
        RECT 22.500 36.280 32.495 36.510 ;
        RECT 33.860 36.280 43.855 36.510 ;
        RECT 23.725 36.250 24.445 36.280 ;
        RECT 41.915 36.270 42.635 36.280 ;
        RECT 22.025 35.920 22.345 36.230 ;
        RECT 31.785 35.870 32.505 35.920 ;
        RECT 32.645 35.900 32.985 36.250 ;
        RECT 33.375 35.900 33.715 36.250 ;
        RECT 33.865 35.870 34.585 35.920 ;
        RECT 44.015 35.890 44.345 36.250 ;
        RECT 22.500 35.640 32.505 35.870 ;
        RECT 33.860 35.640 43.855 35.870 ;
        RECT 31.785 35.600 32.505 35.640 ;
        RECT 33.865 35.590 34.585 35.640 ;
        RECT 22.525 35.310 23.245 35.360 ;
        RECT 33.855 35.310 34.915 35.330 ;
        RECT 43.115 35.310 43.835 35.370 ;
        RECT 22.500 35.080 32.495 35.310 ;
        RECT 33.855 35.080 43.855 35.310 ;
        RECT 22.525 35.040 23.245 35.080 ;
        RECT 33.855 35.070 34.915 35.080 ;
        RECT 43.115 35.030 43.835 35.080 ;
        RECT 22.045 34.970 22.325 35.030 ;
        RECT 21.695 34.780 22.325 34.970 ;
        RECT 21.695 32.570 21.885 34.780 ;
        RECT 22.045 34.720 22.325 34.780 ;
        RECT 32.685 34.720 32.955 35.030 ;
        RECT 33.405 34.720 33.685 35.030 ;
        RECT 44.045 34.970 44.315 35.030 ;
        RECT 44.045 34.780 44.675 34.970 ;
        RECT 44.045 34.720 44.315 34.780 ;
        RECT 31.785 34.670 32.505 34.720 ;
        RECT 33.865 34.670 34.915 34.700 ;
        RECT 22.500 34.440 32.505 34.670 ;
        RECT 33.860 34.440 43.855 34.670 ;
        RECT 31.785 34.400 32.505 34.440 ;
        RECT 33.865 34.390 34.585 34.440 ;
        RECT 23.725 34.110 24.445 34.160 ;
        RECT 41.915 34.110 42.635 34.130 ;
        RECT 22.500 33.880 32.495 34.110 ;
        RECT 33.860 33.880 43.855 34.110 ;
        RECT 23.725 33.850 24.445 33.880 ;
        RECT 41.915 33.870 42.635 33.880 ;
        RECT 22.025 33.520 22.345 33.830 ;
        RECT 31.785 33.470 32.505 33.520 ;
        RECT 32.645 33.500 32.985 33.850 ;
        RECT 33.375 33.500 33.715 33.850 ;
        RECT 33.865 33.470 34.585 33.520 ;
        RECT 44.015 33.490 44.345 33.850 ;
        RECT 22.500 33.240 32.505 33.470 ;
        RECT 33.860 33.240 43.855 33.470 ;
        RECT 31.785 33.200 32.505 33.240 ;
        RECT 33.865 33.190 34.585 33.240 ;
        RECT 22.525 32.910 23.245 32.960 ;
        RECT 33.855 32.910 34.955 32.930 ;
        RECT 43.115 32.910 43.835 32.970 ;
        RECT 22.500 32.680 32.495 32.910 ;
        RECT 33.855 32.680 43.855 32.910 ;
        RECT 22.525 32.640 23.245 32.680 ;
        RECT 33.855 32.670 34.955 32.680 ;
        RECT 43.115 32.630 43.835 32.680 ;
        RECT 22.045 32.570 22.325 32.630 ;
        RECT 21.695 32.380 22.325 32.570 ;
        RECT 22.045 32.320 22.325 32.380 ;
        RECT 32.685 32.320 32.955 32.630 ;
        RECT 33.405 32.320 33.685 32.630 ;
        RECT 44.045 32.570 44.315 32.630 ;
        RECT 44.485 32.570 44.675 34.780 ;
        RECT 44.045 32.380 44.675 32.570 ;
        RECT 44.045 32.320 44.315 32.380 ;
        RECT 31.785 32.270 32.505 32.320 ;
        RECT 33.865 32.270 34.955 32.300 ;
        RECT 22.500 32.040 32.505 32.270 ;
        RECT 33.860 32.040 43.855 32.270 ;
        RECT 31.785 32.000 32.505 32.040 ;
        RECT 33.865 32.030 34.565 32.040 ;
        RECT 44.485 31.390 44.675 32.380 ;
        RECT 18.520 31.130 44.675 31.390 ;
        RECT 28.290 30.060 38.290 30.290 ;
        RECT 28.300 30.030 38.280 30.060 ;
        RECT 27.855 29.950 28.085 30.010 ;
        RECT 38.495 29.950 38.725 30.010 ;
        RECT 27.785 29.110 28.145 29.950 ;
        RECT 38.425 29.110 38.785 29.950 ;
        RECT 27.855 29.050 28.085 29.110 ;
        RECT 38.495 29.050 38.725 29.110 ;
        RECT 28.290 28.770 38.290 29.000 ;
        RECT 7.405 28.520 18.070 28.710 ;
        RECT 29.295 28.690 31.275 28.770 ;
        RECT 35.295 28.690 37.275 28.770 ;
        RECT 7.405 28.480 17.405 28.520 ;
        RECT 6.970 27.470 7.200 28.430 ;
        RECT 17.610 27.790 18.070 28.520 ;
        RECT 19.680 27.790 20.060 27.840 ;
        RECT 17.610 27.530 20.060 27.790 ;
        RECT 17.610 27.470 18.070 27.530 ;
        RECT 19.680 27.490 20.060 27.530 ;
        RECT 20.375 27.790 45.985 28.150 ;
        RECT 7.405 27.190 17.405 27.420 ;
        RECT 7.465 26.930 17.345 27.190 ;
        RECT 6.920 26.850 17.890 26.930 ;
        RECT 6.910 26.620 17.900 26.850 ;
        RECT 20.375 25.560 23.615 27.790 ;
        RECT 23.915 27.170 32.785 27.430 ;
        RECT 34.015 27.420 41.995 27.430 ;
        RECT 34.010 27.190 42.010 27.420 ;
        RECT 34.015 27.170 41.995 27.190 ;
        RECT 23.915 26.780 24.145 27.170 ;
        RECT 32.555 27.080 32.785 27.170 ;
        RECT 33.575 27.080 33.805 27.140 ;
        RECT 32.555 26.780 33.805 27.080 ;
        RECT 42.215 26.780 42.445 27.140 ;
        RECT 23.915 26.520 42.445 26.780 ;
        RECT 23.915 26.180 24.145 26.520 ;
        RECT 32.555 26.240 33.805 26.520 ;
        RECT 32.555 26.180 32.785 26.240 ;
        RECT 33.575 26.180 33.805 26.240 ;
        RECT 42.215 26.180 42.445 26.520 ;
        RECT 24.350 25.900 32.350 26.130 ;
        RECT 34.010 25.900 42.010 26.130 ;
        RECT 24.410 25.560 32.290 25.900 ;
        RECT 34.015 25.560 41.950 25.900 ;
        RECT 42.745 25.560 45.985 27.790 ;
        RECT 6.940 25.260 9.045 25.340 ;
        RECT 15.935 25.330 18.040 25.340 ;
        RECT 6.910 23.500 9.070 25.260 ;
        RECT 15.910 24.390 18.060 25.330 ;
        RECT 20.375 25.290 45.985 25.560 ;
        RECT 20.370 25.180 45.985 25.290 ;
        RECT 20.370 24.910 45.980 25.180 ;
        RECT 15.935 24.030 18.040 24.390 ;
        RECT 19.150 23.500 19.530 23.540 ;
        RECT 6.910 23.240 19.530 23.500 ;
        RECT 1.400 21.030 1.760 22.610 ;
        RECT 6.910 21.450 9.070 23.240 ;
        RECT 19.150 23.190 19.530 23.240 ;
        RECT 15.935 22.710 18.040 22.800 ;
        RECT 1.400 20.770 8.320 21.030 ;
        RECT 1.410 18.900 9.070 20.310 ;
        RECT 15.910 19.345 18.070 22.710 ;
        RECT 20.370 22.680 23.610 24.910 ;
        RECT 24.405 24.570 32.285 24.910 ;
        RECT 34.015 24.570 41.945 24.910 ;
        RECT 24.345 24.340 32.345 24.570 ;
        RECT 34.005 24.340 42.005 24.570 ;
        RECT 23.910 23.950 24.140 24.290 ;
        RECT 32.550 24.230 32.780 24.290 ;
        RECT 33.570 24.230 33.800 24.290 ;
        RECT 32.550 23.950 33.800 24.230 ;
        RECT 42.210 23.950 42.440 24.290 ;
        RECT 23.910 23.690 42.440 23.950 ;
        RECT 23.910 23.300 24.140 23.690 ;
        RECT 32.550 23.390 33.800 23.690 ;
        RECT 32.550 23.300 32.780 23.390 ;
        RECT 33.570 23.330 33.800 23.390 ;
        RECT 42.210 23.330 42.440 23.690 ;
        RECT 23.910 23.040 32.780 23.300 ;
        RECT 34.010 23.280 41.990 23.300 ;
        RECT 34.005 23.050 42.005 23.280 ;
        RECT 34.010 23.040 41.990 23.050 ;
        RECT 42.740 22.680 45.980 24.910 ;
        RECT 20.370 22.320 45.980 22.680 ;
        RECT 29.295 21.700 31.275 21.780 ;
        RECT 35.295 21.700 37.275 21.780 ;
        RECT 28.285 21.470 38.285 21.700 ;
        RECT 27.850 21.360 28.080 21.420 ;
        RECT 38.490 21.360 38.720 21.420 ;
        RECT 27.780 20.520 28.140 21.360 ;
        RECT 38.420 20.520 38.780 21.360 ;
        RECT 27.850 20.460 28.080 20.520 ;
        RECT 38.490 20.460 38.720 20.520 ;
        RECT 28.295 20.410 38.275 20.440 ;
        RECT 28.285 20.180 38.285 20.410 ;
        RECT 15.910 19.340 20.470 19.345 ;
        RECT 15.910 19.080 44.670 19.340 ;
        RECT 15.910 19.075 20.470 19.080 ;
        RECT 15.910 18.900 18.070 19.075 ;
        RECT 1.410 12.410 2.360 18.900 ;
        RECT 25.080 18.640 29.945 18.900 ;
        RECT 19.600 18.370 19.960 18.630 ;
        RECT 31.780 18.430 32.500 18.470 ;
        RECT 33.860 18.430 34.560 18.440 ;
        RECT 6.150 17.560 18.875 17.615 ;
        RECT 2.975 17.530 18.875 17.560 ;
        RECT 2.725 17.525 18.875 17.530 ;
        RECT 2.725 17.360 19.010 17.525 ;
        RECT 2.975 17.355 19.010 17.360 ;
        RECT 2.975 17.330 9.485 17.355 ;
        RECT 3.125 17.090 3.295 17.330 ;
        RECT 3.095 16.090 3.325 17.090 ;
        RECT 3.535 16.080 3.925 17.110 ;
        RECT 4.495 16.970 4.665 16.990 ;
        RECT 6.350 16.970 6.520 17.330 ;
        RECT 8.230 16.970 8.400 17.330 ;
        RECT 9.965 17.325 10.875 17.355 ;
        RECT 11.275 17.325 12.185 17.355 ;
        RECT 12.590 17.325 13.500 17.355 ;
        RECT 13.905 17.325 14.815 17.355 ;
        RECT 15.220 17.325 16.130 17.355 ;
        RECT 16.535 17.325 17.445 17.355 ;
        RECT 17.850 17.325 18.760 17.355 ;
        RECT 10.115 17.085 10.285 17.325 ;
        RECT 3.260 15.900 3.600 15.940 ;
        RECT 3.255 15.640 3.615 15.900 ;
        RECT 3.260 15.600 3.600 15.640 ;
        RECT 3.755 15.290 3.925 16.080 ;
        RECT 4.465 16.260 4.695 16.970 ;
        RECT 5.345 16.260 5.575 16.970 ;
        RECT 4.465 15.680 5.575 16.260 ;
        RECT 3.755 15.120 4.135 15.290 ;
        RECT 3.755 14.625 3.925 15.120 ;
        RECT 4.465 14.970 4.695 15.680 ;
        RECT 5.345 15.100 5.575 15.680 ;
        RECT 5.345 14.950 5.710 15.100 ;
        RECT 6.325 14.970 6.555 16.970 ;
        RECT 7.205 15.100 7.435 16.970 ;
        RECT 7.200 14.950 7.565 15.100 ;
        RECT 8.205 14.970 8.435 16.970 ;
        RECT 9.085 15.100 9.315 16.970 ;
        RECT 10.085 16.085 10.315 17.085 ;
        RECT 10.525 16.075 10.915 17.105 ;
        RECT 11.425 17.085 11.595 17.325 ;
        RECT 11.395 16.085 11.625 17.085 ;
        RECT 11.835 16.075 12.225 17.105 ;
        RECT 12.740 17.085 12.910 17.325 ;
        RECT 12.710 16.085 12.940 17.085 ;
        RECT 13.150 16.075 13.540 17.105 ;
        RECT 14.055 17.085 14.225 17.325 ;
        RECT 14.025 16.085 14.255 17.085 ;
        RECT 14.465 16.075 14.855 17.105 ;
        RECT 15.370 17.085 15.540 17.325 ;
        RECT 15.340 16.085 15.570 17.085 ;
        RECT 15.780 16.075 16.170 17.105 ;
        RECT 16.685 17.085 16.855 17.325 ;
        RECT 16.655 16.085 16.885 17.085 ;
        RECT 17.095 16.075 17.485 17.105 ;
        RECT 18.000 17.085 18.170 17.325 ;
        RECT 17.970 16.085 18.200 17.085 ;
        RECT 18.410 16.075 18.800 17.105 ;
        RECT 10.250 15.895 10.590 15.935 ;
        RECT 10.245 15.635 10.605 15.895 ;
        RECT 10.250 15.595 10.590 15.635 ;
        RECT 10.745 15.285 10.915 16.075 ;
        RECT 11.560 15.895 11.900 15.935 ;
        RECT 11.555 15.635 11.915 15.895 ;
        RECT 11.560 15.595 11.900 15.635 ;
        RECT 11.645 15.330 11.815 15.595 ;
        RECT 11.645 15.285 11.810 15.330 ;
        RECT 10.745 15.115 11.810 15.285 ;
        RECT 12.055 15.285 12.225 16.075 ;
        RECT 12.875 15.895 13.215 15.935 ;
        RECT 12.870 15.635 13.230 15.895 ;
        RECT 12.875 15.595 13.215 15.635 ;
        RECT 13.370 15.285 13.540 16.075 ;
        RECT 14.190 15.895 14.530 15.935 ;
        RECT 14.185 15.635 14.545 15.895 ;
        RECT 14.190 15.595 14.530 15.635 ;
        RECT 14.270 15.285 14.440 15.595 ;
        RECT 12.055 15.115 14.440 15.285 ;
        RECT 14.685 15.285 14.855 16.075 ;
        RECT 15.505 15.895 15.845 15.935 ;
        RECT 15.500 15.635 15.860 15.895 ;
        RECT 15.505 15.595 15.845 15.635 ;
        RECT 16.000 15.285 16.170 16.075 ;
        RECT 16.820 15.895 17.160 15.935 ;
        RECT 16.815 15.635 17.175 15.895 ;
        RECT 16.820 15.595 17.160 15.635 ;
        RECT 17.315 15.285 17.485 16.075 ;
        RECT 18.135 15.895 18.475 15.935 ;
        RECT 18.130 15.635 18.490 15.895 ;
        RECT 18.135 15.595 18.475 15.635 ;
        RECT 18.630 15.285 18.800 16.075 ;
        RECT 14.685 15.115 19.230 15.285 ;
        RECT 9.080 14.950 9.445 15.100 ;
        RECT 4.535 14.625 4.865 14.705 ;
        RECT 3.755 14.455 4.865 14.625 ;
        RECT 3.260 14.230 3.595 14.270 ;
        RECT 3.245 13.970 3.605 14.230 ;
        RECT 3.260 13.930 3.595 13.970 ;
        RECT 3.755 13.750 3.925 14.455 ;
        RECT 4.535 14.375 4.865 14.455 ;
        RECT 4.165 14.205 4.525 14.230 ;
        RECT 5.080 14.205 5.420 14.290 ;
        RECT 4.100 14.035 5.420 14.205 ;
        RECT 4.165 13.960 4.525 14.035 ;
        RECT 5.080 13.950 5.420 14.035 ;
        RECT 5.560 13.840 5.710 14.950 ;
        RECT 6.475 14.780 6.815 14.820 ;
        RECT 6.465 14.735 6.825 14.780 ;
        RECT 5.955 14.565 6.825 14.735 ;
        RECT 6.465 14.520 6.825 14.565 ;
        RECT 7.415 14.735 7.565 14.950 ;
        RECT 8.355 14.735 8.695 14.820 ;
        RECT 7.415 14.565 8.695 14.735 ;
        RECT 6.475 14.480 6.815 14.520 ;
        RECT 6.935 14.260 7.275 14.290 ;
        RECT 6.885 14.205 7.275 14.260 ;
        RECT 5.955 14.035 7.275 14.205 ;
        RECT 6.885 14.000 7.275 14.035 ;
        RECT 6.935 13.950 7.275 14.000 ;
        RECT 5.560 13.770 6.165 13.840 ;
        RECT 7.415 13.770 7.565 14.565 ;
        RECT 8.355 14.480 8.695 14.565 ;
        RECT 9.295 14.780 9.445 14.950 ;
        RECT 9.295 14.520 9.715 14.780 ;
        RECT 7.745 14.205 8.105 14.250 ;
        RECT 8.815 14.205 9.155 14.290 ;
        RECT 7.745 14.035 9.155 14.205 ;
        RECT 7.745 13.990 8.105 14.035 ;
        RECT 8.815 13.950 9.155 14.035 ;
        RECT 9.295 13.770 9.445 14.520 ;
        RECT 10.250 14.225 10.585 14.265 ;
        RECT 10.235 13.965 10.595 14.225 ;
        RECT 10.250 13.925 10.585 13.965 ;
        RECT 3.095 12.750 3.325 13.750 ;
        RECT 3.125 12.510 3.295 12.750 ;
        RECT 3.535 12.730 3.925 13.750 ;
        RECT 4.465 12.750 4.695 13.750 ;
        RECT 5.345 13.620 6.165 13.770 ;
        RECT 6.350 13.750 7.565 13.770 ;
        RECT 8.230 13.750 9.445 13.770 ;
        RECT 4.495 12.510 4.665 12.750 ;
        RECT 5.345 12.745 5.575 13.620 ;
        RECT 5.805 13.580 6.165 13.620 ;
        RECT 6.320 13.620 7.565 13.750 ;
        RECT 8.200 13.620 9.445 13.750 ;
        RECT 10.745 13.745 10.915 15.115 ;
        RECT 11.560 14.225 11.895 14.265 ;
        RECT 11.545 13.965 11.905 14.225 ;
        RECT 11.560 13.925 11.895 13.965 ;
        RECT 12.055 13.745 12.225 15.115 ;
        RECT 12.875 14.225 13.210 14.265 ;
        RECT 12.860 13.965 13.220 14.225 ;
        RECT 12.875 13.925 13.210 13.965 ;
        RECT 13.370 13.745 13.540 15.115 ;
        RECT 14.190 14.225 14.525 14.265 ;
        RECT 14.175 13.965 14.535 14.225 ;
        RECT 14.190 13.925 14.525 13.965 ;
        RECT 14.685 13.745 14.855 15.115 ;
        RECT 15.505 14.225 15.840 14.265 ;
        RECT 15.490 13.965 15.850 14.225 ;
        RECT 15.505 13.925 15.840 13.965 ;
        RECT 16.000 13.745 16.170 15.115 ;
        RECT 16.820 14.225 17.155 14.265 ;
        RECT 16.805 13.965 17.165 14.225 ;
        RECT 16.820 13.925 17.155 13.965 ;
        RECT 17.315 13.745 17.485 15.115 ;
        RECT 18.135 14.225 18.470 14.265 ;
        RECT 18.120 13.965 18.480 14.225 ;
        RECT 18.135 13.925 18.470 13.965 ;
        RECT 18.630 13.745 18.800 15.115 ;
        RECT 6.320 12.750 6.550 13.620 ;
        RECT 7.200 13.160 7.430 13.620 ;
        RECT 7.135 12.900 7.495 13.160 ;
        RECT 7.200 12.745 7.430 12.900 ;
        RECT 8.200 12.750 8.430 13.620 ;
        RECT 9.080 12.745 9.310 13.620 ;
        RECT 10.085 12.745 10.315 13.745 ;
        RECT 2.975 12.480 3.885 12.510 ;
        RECT 4.345 12.480 5.695 12.510 ;
        RECT 6.200 12.480 7.550 12.510 ;
        RECT 8.080 12.480 9.430 12.510 ;
        RECT 10.115 12.505 10.285 12.745 ;
        RECT 10.525 12.740 10.915 13.745 ;
        RECT 11.395 12.745 11.625 13.745 ;
        RECT 10.555 12.725 10.915 12.740 ;
        RECT 11.425 12.505 11.595 12.745 ;
        RECT 11.835 12.740 12.225 13.745 ;
        RECT 12.710 12.745 12.940 13.745 ;
        RECT 11.865 12.725 12.225 12.740 ;
        RECT 12.740 12.505 12.910 12.745 ;
        RECT 13.150 12.740 13.540 13.745 ;
        RECT 14.025 12.745 14.255 13.745 ;
        RECT 13.180 12.725 13.540 12.740 ;
        RECT 14.055 12.505 14.225 12.745 ;
        RECT 14.465 12.740 14.855 13.745 ;
        RECT 15.340 12.745 15.570 13.745 ;
        RECT 14.495 12.725 14.855 12.740 ;
        RECT 15.370 12.505 15.540 12.745 ;
        RECT 15.780 12.740 16.170 13.745 ;
        RECT 16.655 12.745 16.885 13.745 ;
        RECT 15.810 12.725 16.170 12.740 ;
        RECT 16.685 12.505 16.855 12.745 ;
        RECT 17.095 12.740 17.485 13.745 ;
        RECT 17.970 12.745 18.200 13.745 ;
        RECT 17.125 12.725 17.485 12.740 ;
        RECT 18.000 12.505 18.170 12.745 ;
        RECT 18.410 12.740 18.800 13.745 ;
        RECT 18.440 12.725 18.800 12.740 ;
        RECT 2.975 12.410 3.905 12.480 ;
        RECT 4.305 12.475 9.430 12.480 ;
        RECT 9.965 12.475 10.875 12.505 ;
        RECT 11.275 12.475 12.185 12.505 ;
        RECT 12.590 12.475 13.500 12.505 ;
        RECT 13.905 12.475 14.815 12.505 ;
        RECT 15.220 12.475 16.130 12.505 ;
        RECT 16.535 12.475 17.445 12.505 ;
        RECT 17.850 12.475 18.760 12.505 ;
        RECT 4.305 12.410 18.760 12.475 ;
        RECT 1.410 12.275 18.760 12.410 ;
        RECT 1.410 11.730 18.700 12.275 ;
        RECT 1.410 11.700 17.810 11.730 ;
        RECT 1.410 7.640 6.690 11.700 ;
        RECT 7.570 11.360 10.500 11.420 ;
        RECT 7.360 11.130 17.360 11.360 ;
        RECT 6.970 8.190 7.200 11.100 ;
        RECT 17.520 11.020 17.750 11.100 ;
        RECT 19.060 11.020 19.230 15.115 ;
        RECT 19.650 13.390 19.910 18.370 ;
        RECT 22.495 18.200 32.500 18.430 ;
        RECT 33.855 18.200 43.850 18.430 ;
        RECT 31.780 18.150 32.500 18.200 ;
        RECT 33.860 18.170 34.950 18.200 ;
        RECT 22.040 18.090 22.320 18.150 ;
        RECT 21.690 17.900 22.320 18.090 ;
        RECT 21.690 15.690 21.880 17.900 ;
        RECT 22.040 17.840 22.320 17.900 ;
        RECT 32.680 17.840 32.950 18.150 ;
        RECT 33.400 17.840 33.680 18.150 ;
        RECT 44.040 18.090 44.310 18.150 ;
        RECT 44.480 18.090 44.670 19.080 ;
        RECT 44.040 17.900 44.670 18.090 ;
        RECT 44.040 17.840 44.310 17.900 ;
        RECT 22.520 17.790 23.240 17.830 ;
        RECT 33.850 17.790 34.950 17.800 ;
        RECT 43.110 17.790 43.830 17.840 ;
        RECT 22.495 17.560 32.490 17.790 ;
        RECT 33.850 17.560 43.850 17.790 ;
        RECT 22.520 17.510 23.240 17.560 ;
        RECT 33.850 17.540 34.950 17.560 ;
        RECT 43.110 17.500 43.830 17.560 ;
        RECT 31.780 17.230 32.500 17.270 ;
        RECT 33.860 17.230 34.580 17.280 ;
        RECT 22.495 17.000 32.500 17.230 ;
        RECT 33.855 17.000 43.850 17.230 ;
        RECT 31.780 16.950 32.500 17.000 ;
        RECT 22.020 16.640 22.340 16.950 ;
        RECT 32.640 16.620 32.980 16.970 ;
        RECT 33.370 16.620 33.710 16.970 ;
        RECT 33.860 16.950 34.580 17.000 ;
        RECT 44.010 16.620 44.340 16.980 ;
        RECT 23.720 16.590 24.440 16.620 ;
        RECT 41.910 16.590 42.630 16.600 ;
        RECT 22.495 16.360 32.490 16.590 ;
        RECT 33.855 16.360 43.850 16.590 ;
        RECT 23.720 16.310 24.440 16.360 ;
        RECT 41.910 16.340 42.630 16.360 ;
        RECT 31.780 16.030 32.500 16.070 ;
        RECT 33.860 16.030 34.580 16.080 ;
        RECT 22.495 15.800 32.500 16.030 ;
        RECT 33.855 15.800 43.850 16.030 ;
        RECT 31.780 15.750 32.500 15.800 ;
        RECT 33.860 15.770 34.910 15.800 ;
        RECT 22.040 15.690 22.320 15.750 ;
        RECT 21.690 15.500 22.320 15.690 ;
        RECT 21.690 13.390 21.880 15.500 ;
        RECT 22.040 15.440 22.320 15.500 ;
        RECT 32.680 15.440 32.950 15.750 ;
        RECT 33.400 15.440 33.680 15.750 ;
        RECT 44.040 15.690 44.310 15.750 ;
        RECT 44.480 15.690 44.670 17.900 ;
        RECT 44.040 15.500 44.670 15.690 ;
        RECT 44.040 15.440 44.310 15.500 ;
        RECT 22.520 15.390 23.240 15.430 ;
        RECT 33.850 15.390 34.910 15.400 ;
        RECT 43.110 15.390 43.830 15.440 ;
        RECT 22.495 15.160 32.490 15.390 ;
        RECT 33.850 15.160 43.850 15.390 ;
        RECT 22.520 15.110 23.240 15.160 ;
        RECT 33.850 15.140 34.910 15.160 ;
        RECT 43.110 15.100 43.830 15.160 ;
        RECT 31.780 14.830 32.500 14.870 ;
        RECT 33.860 14.830 34.580 14.880 ;
        RECT 22.495 14.600 32.500 14.830 ;
        RECT 33.855 14.600 43.850 14.830 ;
        RECT 31.780 14.550 32.500 14.600 ;
        RECT 22.020 14.240 22.340 14.550 ;
        RECT 32.640 14.220 32.980 14.570 ;
        RECT 33.370 14.220 33.710 14.570 ;
        RECT 33.860 14.550 34.580 14.600 ;
        RECT 44.010 14.220 44.340 14.580 ;
        RECT 23.720 14.190 24.440 14.220 ;
        RECT 41.910 14.190 42.630 14.200 ;
        RECT 22.495 13.960 32.490 14.190 ;
        RECT 33.855 13.960 43.850 14.190 ;
        RECT 23.720 13.910 24.440 13.960 ;
        RECT 41.910 13.940 42.630 13.960 ;
        RECT 19.650 13.130 44.340 13.390 ;
        RECT 23.710 12.730 43.830 12.990 ;
        RECT 22.510 12.330 42.630 12.590 ;
        RECT 17.520 10.830 19.230 11.020 ;
        RECT 21.030 11.450 25.410 11.470 ;
        RECT 27.280 11.450 32.260 11.470 ;
        RECT 34.250 11.450 39.230 11.470 ;
        RECT 21.030 11.210 25.810 11.450 ;
        RECT 27.270 11.220 32.270 11.450 ;
        RECT 34.240 11.220 39.240 11.450 ;
        RECT 27.280 11.210 32.260 11.220 ;
        RECT 34.250 11.210 39.230 11.220 ;
        RECT 40.570 11.210 45.320 11.470 ;
        RECT 14.290 10.720 17.220 10.780 ;
        RECT 7.360 10.490 17.360 10.720 ;
        RECT 7.570 10.080 10.500 10.140 ;
        RECT 7.360 9.850 17.360 10.080 ;
        RECT 14.290 9.440 17.220 9.500 ;
        RECT 7.360 9.210 17.360 9.440 ;
        RECT 7.570 8.800 10.500 8.860 ;
        RECT 7.360 8.570 17.360 8.800 ;
        RECT 17.520 8.190 17.750 10.830 ;
        RECT 21.030 10.820 21.260 11.210 ;
        RECT 25.580 11.110 25.810 11.210 ;
        RECT 40.570 11.190 40.930 11.210 ;
        RECT 40.570 11.170 40.770 11.190 ;
        RECT 26.880 11.110 27.110 11.170 ;
        RECT 32.430 11.110 32.660 11.170 ;
        RECT 33.850 11.110 34.080 11.170 ;
        RECT 39.400 11.110 39.630 11.170 ;
        RECT 40.540 11.110 40.770 11.170 ;
        RECT 25.580 10.820 27.110 11.110 ;
        RECT 32.360 10.820 32.720 11.110 ;
        RECT 21.030 10.560 32.720 10.820 ;
        RECT 21.030 10.210 21.260 10.560 ;
        RECT 25.580 10.270 27.110 10.560 ;
        RECT 32.360 10.270 32.720 10.560 ;
        RECT 33.790 10.820 34.150 11.110 ;
        RECT 39.400 10.820 40.770 11.110 ;
        RECT 45.090 10.820 45.320 11.210 ;
        RECT 33.790 10.560 45.320 10.820 ;
        RECT 33.790 10.270 34.150 10.560 ;
        RECT 39.400 10.270 40.770 10.560 ;
        RECT 25.580 10.210 25.810 10.270 ;
        RECT 26.880 10.210 27.110 10.270 ;
        RECT 32.430 10.210 32.660 10.270 ;
        RECT 33.850 10.210 34.080 10.270 ;
        RECT 39.400 10.210 39.630 10.270 ;
        RECT 40.540 10.210 40.770 10.270 ;
        RECT 45.090 10.210 45.320 10.560 ;
        RECT 21.420 9.930 25.420 10.160 ;
        RECT 27.270 9.930 32.270 10.160 ;
        RECT 34.240 9.930 39.240 10.160 ;
        RECT 40.930 9.930 44.930 10.160 ;
        RECT 21.730 9.560 25.100 9.930 ;
        RECT 28.020 9.560 31.390 9.930 ;
        RECT 35.130 9.560 38.500 9.930 ;
        RECT 20.370 9.390 45.980 9.560 ;
        RECT 7.360 7.930 17.360 8.160 ;
        RECT 14.290 7.870 17.220 7.930 ;
        RECT 20.370 7.640 26.290 9.390 ;
        RECT 27.280 9.020 32.260 9.040 ;
        RECT 34.250 9.020 39.230 9.040 ;
        RECT 27.270 8.790 32.270 9.020 ;
        RECT 34.240 8.790 39.240 9.020 ;
        RECT 27.280 8.780 32.260 8.790 ;
        RECT 34.250 8.780 39.230 8.790 ;
        RECT 26.880 8.400 27.110 8.740 ;
        RECT 32.430 8.680 32.660 8.740 ;
        RECT 33.850 8.680 34.080 8.740 ;
        RECT 32.360 8.400 32.720 8.680 ;
        RECT 26.880 8.140 32.720 8.400 ;
        RECT 26.880 7.780 27.110 8.140 ;
        RECT 32.360 7.840 32.720 8.140 ;
        RECT 33.790 8.400 34.150 8.680 ;
        RECT 39.400 8.400 39.630 8.740 ;
        RECT 33.790 8.140 39.630 8.400 ;
        RECT 33.790 7.840 34.150 8.140 ;
        RECT 32.430 7.780 32.660 7.840 ;
        RECT 33.850 7.780 34.080 7.840 ;
        RECT 39.400 7.780 39.630 8.140 ;
        RECT 27.270 7.640 32.270 7.730 ;
        RECT 34.240 7.640 39.240 7.730 ;
        RECT 40.060 7.640 45.980 9.390 ;
        RECT 1.410 7.330 45.980 7.640 ;
        RECT 1.410 7.130 45.990 7.330 ;
        RECT 1.410 5.130 46.035 7.130 ;
        RECT 7.570 1.430 13.540 2.150 ;
      LAYER via ;
        RECT 5.230 50.840 5.500 52.070 ;
        RECT 7.110 50.940 7.380 52.170 ;
        RECT 18.520 46.690 20.530 46.950 ;
        RECT 12.630 42.330 17.510 42.610 ;
        RECT 22.100 45.740 24.110 46.000 ;
        RECT 20.545 43.340 45.805 43.620 ;
        RECT 19.570 41.610 19.830 41.870 ;
        RECT 32.415 41.790 32.675 42.630 ;
        RECT 33.845 41.790 34.105 42.630 ;
        RECT 27.335 41.430 32.215 41.690 ;
        RECT 34.305 41.430 39.185 41.690 ;
        RECT 32.415 39.360 32.675 40.200 ;
        RECT 33.845 39.360 34.105 40.200 ;
        RECT 21.485 39.000 25.365 39.260 ;
        RECT 27.335 39.000 32.215 39.260 ;
        RECT 34.305 39.000 39.185 39.260 ;
        RECT 40.985 39.000 44.865 39.260 ;
        RECT 22.565 37.880 23.195 38.140 ;
        RECT 41.955 37.880 42.585 38.140 ;
        RECT 23.765 37.480 24.395 37.740 ;
        RECT 43.165 37.480 43.795 37.740 ;
        RECT 19.180 37.070 19.500 37.360 ;
        RECT 33.415 37.080 33.675 37.340 ;
        RECT 44.055 37.080 44.315 37.340 ;
        RECT 23.765 36.270 24.395 36.530 ;
        RECT 41.965 36.270 42.595 36.530 ;
        RECT 22.055 35.940 22.315 36.200 ;
        RECT 32.685 35.950 32.945 36.210 ;
        RECT 33.425 35.950 33.685 36.210 ;
        RECT 44.045 35.940 44.305 36.200 ;
        RECT 31.825 35.630 32.455 35.890 ;
        RECT 33.905 35.630 34.535 35.890 ;
        RECT 22.565 35.070 23.195 35.330 ;
        RECT 43.165 35.070 43.795 35.330 ;
        RECT 31.825 34.430 32.455 34.690 ;
        RECT 33.905 34.430 34.535 34.690 ;
        RECT 23.765 33.870 24.395 34.130 ;
        RECT 41.965 33.870 42.595 34.130 ;
        RECT 22.055 33.540 22.315 33.800 ;
        RECT 32.685 33.550 32.945 33.810 ;
        RECT 33.425 33.550 33.685 33.810 ;
        RECT 44.045 33.540 44.305 33.800 ;
        RECT 31.825 33.230 32.455 33.490 ;
        RECT 33.905 33.230 34.535 33.490 ;
        RECT 22.565 32.670 23.195 32.930 ;
        RECT 43.165 32.670 43.795 32.930 ;
        RECT 31.825 32.030 32.455 32.290 ;
        RECT 33.905 32.030 34.535 32.290 ;
        RECT 22.055 31.130 22.315 31.390 ;
        RECT 32.685 31.130 32.945 31.390 ;
        RECT 28.350 30.030 38.230 30.290 ;
        RECT 27.835 29.110 28.095 29.950 ;
        RECT 38.475 29.110 38.735 29.950 ;
        RECT 29.345 28.690 31.225 28.970 ;
        RECT 35.345 28.690 37.225 28.970 ;
        RECT 19.710 27.520 20.030 27.810 ;
        RECT 6.970 26.650 17.840 26.930 ;
        RECT 24.405 27.170 32.285 27.430 ;
        RECT 34.065 27.170 41.945 27.430 ;
        RECT 15.960 24.390 18.010 25.330 ;
        RECT 1.450 20.770 1.710 22.610 ;
        RECT 19.180 23.220 19.500 23.510 ;
        RECT 8.010 20.770 8.270 21.030 ;
        RECT 34.065 24.375 36.870 26.100 ;
        RECT 24.400 23.040 32.280 23.300 ;
        RECT 34.060 23.040 41.940 23.300 ;
        RECT 29.345 21.500 31.225 21.780 ;
        RECT 35.345 21.500 37.225 21.780 ;
        RECT 27.830 20.520 28.090 21.360 ;
        RECT 38.470 20.520 38.730 21.360 ;
        RECT 28.345 20.180 38.225 20.440 ;
        RECT 22.050 19.080 22.310 19.340 ;
        RECT 32.680 19.080 32.940 19.340 ;
        RECT 25.130 18.640 29.895 18.900 ;
        RECT 19.650 18.370 19.910 18.630 ;
        RECT 6.200 17.355 18.825 17.615 ;
        RECT 3.305 15.640 3.565 15.900 ;
        RECT 10.295 15.635 10.555 15.895 ;
        RECT 11.605 15.635 11.865 15.895 ;
        RECT 12.920 15.635 13.180 15.895 ;
        RECT 14.235 15.635 14.495 15.895 ;
        RECT 15.550 15.635 15.810 15.895 ;
        RECT 16.865 15.635 17.125 15.895 ;
        RECT 18.180 15.635 18.440 15.895 ;
        RECT 3.295 13.970 3.555 14.230 ;
        RECT 4.215 13.960 4.475 14.230 ;
        RECT 6.515 14.520 6.775 14.780 ;
        RECT 6.935 14.000 7.195 14.260 ;
        RECT 5.855 13.580 6.115 13.840 ;
        RECT 9.405 14.520 9.665 14.780 ;
        RECT 7.795 13.990 8.055 14.250 ;
        RECT 10.285 13.965 10.545 14.225 ;
        RECT 11.595 13.965 11.855 14.225 ;
        RECT 12.910 13.965 13.170 14.225 ;
        RECT 14.225 13.965 14.485 14.225 ;
        RECT 15.540 13.965 15.800 14.225 ;
        RECT 16.855 13.965 17.115 14.225 ;
        RECT 18.170 13.965 18.430 14.225 ;
        RECT 7.185 12.900 7.445 13.160 ;
        RECT 7.620 11.160 10.450 11.420 ;
        RECT 31.820 18.180 32.450 18.440 ;
        RECT 33.900 18.180 34.530 18.440 ;
        RECT 22.560 17.540 23.190 17.800 ;
        RECT 43.160 17.540 43.790 17.800 ;
        RECT 31.820 16.980 32.450 17.240 ;
        RECT 33.900 16.980 34.530 17.240 ;
        RECT 22.050 16.670 22.310 16.930 ;
        RECT 32.680 16.660 32.940 16.920 ;
        RECT 33.420 16.660 33.680 16.920 ;
        RECT 44.040 16.670 44.300 16.930 ;
        RECT 23.760 16.340 24.390 16.600 ;
        RECT 41.960 16.340 42.590 16.600 ;
        RECT 31.820 15.780 32.450 16.040 ;
        RECT 33.900 15.780 34.530 16.040 ;
        RECT 22.560 15.140 23.190 15.400 ;
        RECT 43.160 15.140 43.790 15.400 ;
        RECT 31.820 14.580 32.450 14.840 ;
        RECT 33.900 14.580 34.530 14.840 ;
        RECT 22.050 14.270 22.310 14.530 ;
        RECT 32.680 14.260 32.940 14.520 ;
        RECT 33.420 14.260 33.680 14.520 ;
        RECT 44.040 14.270 44.300 14.530 ;
        RECT 23.760 13.940 24.390 14.200 ;
        RECT 41.960 13.940 42.590 14.200 ;
        RECT 33.410 13.130 33.670 13.390 ;
        RECT 44.050 13.130 44.310 13.390 ;
        RECT 23.760 12.730 24.390 12.990 ;
        RECT 43.160 12.730 43.790 12.990 ;
        RECT 22.560 12.330 23.190 12.590 ;
        RECT 41.950 12.330 42.580 12.590 ;
        RECT 21.480 11.210 25.360 11.470 ;
        RECT 27.330 11.210 32.210 11.470 ;
        RECT 34.300 11.210 39.180 11.470 ;
        RECT 40.980 11.210 44.860 11.470 ;
        RECT 14.340 10.520 17.170 10.780 ;
        RECT 7.620 9.880 10.450 10.140 ;
        RECT 14.340 9.240 17.170 9.500 ;
        RECT 7.620 8.600 10.450 8.860 ;
        RECT 32.410 10.270 32.670 11.110 ;
        RECT 33.840 10.270 34.100 11.110 ;
        RECT 14.340 7.870 17.170 8.130 ;
        RECT 27.330 8.780 32.210 9.040 ;
        RECT 34.300 8.780 39.180 9.040 ;
        RECT 32.410 7.840 32.670 8.680 ;
        RECT 33.840 7.840 34.100 8.680 ;
        RECT 14.420 7.330 17.070 7.610 ;
        RECT 20.540 6.850 45.800 7.130 ;
        RECT 7.620 1.430 13.490 2.150 ;
      LAYER met2 ;
        RECT 5.180 50.790 5.550 52.120 ;
        RECT 7.060 50.890 7.430 52.220 ;
        RECT 5.235 50.085 5.505 50.790 ;
        RECT 1.440 49.815 5.505 50.085 ;
        RECT 1.440 45.370 1.710 49.815 ;
        RECT 7.115 48.695 7.385 50.890 ;
        RECT 1.880 48.425 7.385 48.695 ;
        RECT 1.880 45.395 2.150 48.425 ;
        RECT 18.520 46.590 20.530 47.050 ;
        RECT 22.100 45.640 24.110 46.100 ;
        RECT 1.450 20.720 1.710 45.370 ;
        RECT 1.850 12.730 2.170 45.395 ;
        RECT 20.545 43.290 45.805 43.670 ;
        RECT 2.315 42.890 45.860 43.150 ;
        RECT 2.315 15.910 2.575 42.890 ;
        RECT 12.630 42.280 17.510 42.660 ;
        RECT 19.570 40.590 19.830 41.920 ;
        RECT 27.335 41.690 32.215 41.740 ;
        RECT 18.560 40.330 19.830 40.590 ;
        RECT 20.505 41.430 32.215 41.690 ;
        RECT 6.970 26.600 17.840 26.980 ;
        RECT 15.960 24.340 18.010 25.380 ;
        RECT 18.560 22.030 18.820 40.330 ;
        RECT 19.150 37.040 19.530 37.390 ;
        RECT 19.210 23.540 19.470 37.040 ;
        RECT 19.680 27.490 20.060 27.840 ;
        RECT 19.740 25.870 20.000 27.490 ;
        RECT 20.505 27.430 20.765 41.430 ;
        RECT 27.335 41.380 32.215 41.430 ;
        RECT 32.415 39.310 32.675 42.680 ;
        RECT 33.845 39.310 34.105 42.680 ;
        RECT 34.305 41.690 39.185 41.740 ;
        RECT 45.600 41.690 45.860 42.890 ;
        RECT 34.305 41.580 45.860 41.690 ;
        RECT 34.305 41.430 45.855 41.580 ;
        RECT 34.305 41.380 39.185 41.430 ;
        RECT 21.485 38.950 25.365 39.310 ;
        RECT 27.335 38.950 32.215 39.310 ;
        RECT 34.305 38.950 39.185 39.310 ;
        RECT 40.985 38.950 44.865 39.310 ;
        RECT 22.015 35.900 22.355 36.250 ;
        RECT 22.015 33.850 22.345 35.900 ;
        RECT 22.015 31.130 22.355 33.850 ;
        RECT 22.525 32.640 23.245 38.950 ;
        RECT 27.335 38.790 27.595 38.950 ;
        RECT 24.185 38.530 27.595 38.790 ;
        RECT 38.925 38.790 39.185 38.950 ;
        RECT 38.925 38.530 42.175 38.790 ;
        RECT 24.185 37.810 24.445 38.530 ;
        RECT 27.335 38.520 27.595 38.530 ;
        RECT 23.725 33.850 24.445 37.810 ;
        RECT 41.915 38.190 42.175 38.530 ;
        RECT 41.915 38.140 42.585 38.190 ;
        RECT 31.785 30.825 32.505 35.900 ;
        RECT 32.645 31.130 32.985 36.250 ;
        RECT 33.375 33.500 33.715 37.340 ;
        RECT 33.865 30.825 34.585 35.920 ;
        RECT 41.915 33.870 42.635 38.140 ;
        RECT 43.115 32.630 43.835 38.950 ;
        RECT 44.015 33.490 44.345 37.340 ;
        RECT 31.775 30.340 34.585 30.825 ;
        RECT 27.835 29.660 28.095 30.000 ;
        RECT 28.350 29.980 38.230 30.340 ;
        RECT 33.045 29.660 33.305 29.670 ;
        RECT 38.475 29.660 38.735 30.000 ;
        RECT 27.835 29.400 38.735 29.660 ;
        RECT 27.835 29.060 28.095 29.400 ;
        RECT 29.345 28.640 31.225 29.020 ;
        RECT 24.405 27.430 32.285 27.480 ;
        RECT 20.505 27.170 32.285 27.430 ;
        RECT 24.405 27.120 32.285 27.170 ;
        RECT 33.045 25.870 33.305 29.400 ;
        RECT 38.475 29.060 38.735 29.400 ;
        RECT 35.345 28.640 37.225 29.020 ;
        RECT 34.065 27.430 41.945 27.480 ;
        RECT 45.595 27.430 45.855 41.430 ;
        RECT 34.065 27.170 45.985 27.430 ;
        RECT 34.065 27.120 41.945 27.170 ;
        RECT 19.740 25.610 33.305 25.870 ;
        RECT 19.740 24.860 20.000 25.610 ;
        RECT 19.740 24.600 33.300 24.860 ;
        RECT 19.150 23.190 19.530 23.540 ;
        RECT 24.400 23.300 32.280 23.350 ;
        RECT 20.500 23.040 32.280 23.300 ;
        RECT 18.560 21.770 19.910 22.030 ;
        RECT 8.010 21.030 8.270 21.080 ;
        RECT 8.010 20.770 19.370 21.030 ;
        RECT 8.010 20.720 8.270 20.770 ;
        RECT 6.200 17.305 18.825 17.685 ;
        RECT 2.725 17.065 4.120 17.245 ;
        RECT 2.725 17.060 3.145 17.065 ;
        RECT 3.305 15.940 3.565 15.950 ;
        RECT 2.985 15.910 3.605 15.940 ;
        RECT 2.315 15.640 3.605 15.910 ;
        RECT 2.725 15.630 3.605 15.640 ;
        RECT 2.985 15.600 3.605 15.630 ;
        RECT 3.305 15.590 3.565 15.600 ;
        RECT 3.345 14.280 3.515 15.590 ;
        RECT 3.950 14.795 4.120 17.065 ;
        RECT 10.295 15.935 10.555 15.945 ;
        RECT 11.605 15.935 11.865 15.945 ;
        RECT 12.920 15.935 13.180 15.945 ;
        RECT 14.235 15.935 14.495 15.945 ;
        RECT 15.550 15.935 15.810 15.945 ;
        RECT 16.865 15.935 17.125 15.945 ;
        RECT 18.180 15.935 18.440 15.945 ;
        RECT 9.715 15.895 9.985 15.905 ;
        RECT 9.700 15.850 9.985 15.895 ;
        RECT 10.245 15.850 10.595 15.935 ;
        RECT 9.700 15.680 10.595 15.850 ;
        RECT 9.700 15.625 9.985 15.680 ;
        RECT 9.700 14.830 9.870 15.625 ;
        RECT 10.245 15.595 10.595 15.680 ;
        RECT 11.025 15.850 11.295 15.905 ;
        RECT 11.555 15.850 11.905 15.935 ;
        RECT 12.340 15.850 12.610 15.905 ;
        RECT 12.870 15.850 13.220 15.935 ;
        RECT 11.025 15.680 13.220 15.850 ;
        RECT 11.025 15.625 11.295 15.680 ;
        RECT 11.555 15.595 11.905 15.680 ;
        RECT 12.340 15.625 12.610 15.680 ;
        RECT 12.870 15.595 13.220 15.680 ;
        RECT 13.655 15.850 13.925 15.905 ;
        RECT 14.185 15.850 14.535 15.935 ;
        RECT 14.970 15.850 15.240 15.905 ;
        RECT 15.500 15.850 15.850 15.935 ;
        RECT 16.285 15.850 16.555 15.905 ;
        RECT 16.815 15.850 17.165 15.935 ;
        RECT 17.600 15.850 17.870 15.905 ;
        RECT 18.130 15.895 18.480 15.935 ;
        RECT 19.110 15.895 19.370 20.770 ;
        RECT 19.650 18.320 19.910 21.770 ;
        RECT 18.130 15.850 19.370 15.895 ;
        RECT 13.655 15.680 19.370 15.850 ;
        RECT 13.655 15.625 13.925 15.680 ;
        RECT 14.185 15.595 14.535 15.680 ;
        RECT 14.970 15.625 15.240 15.680 ;
        RECT 15.500 15.595 15.850 15.680 ;
        RECT 16.285 15.625 16.555 15.680 ;
        RECT 16.815 15.595 17.165 15.680 ;
        RECT 17.600 15.625 17.870 15.680 ;
        RECT 18.130 15.635 19.370 15.680 ;
        RECT 18.130 15.595 18.480 15.635 ;
        RECT 19.110 15.630 19.370 15.635 ;
        RECT 10.295 15.585 10.555 15.595 ;
        RECT 11.605 15.585 11.865 15.595 ;
        RECT 12.920 15.585 13.180 15.595 ;
        RECT 14.235 15.585 14.495 15.595 ;
        RECT 15.550 15.585 15.810 15.595 ;
        RECT 16.865 15.585 17.125 15.595 ;
        RECT 18.180 15.585 18.440 15.595 ;
        RECT 3.950 14.625 5.590 14.795 ;
        RECT 3.295 13.920 3.555 14.280 ;
        RECT 4.215 13.660 4.475 14.280 ;
        RECT 5.320 14.205 5.590 14.625 ;
        RECT 6.515 14.735 6.775 14.830 ;
        RECT 9.405 14.735 9.870 14.830 ;
        RECT 6.515 14.565 9.870 14.735 ;
        RECT 6.515 14.470 6.775 14.565 ;
        RECT 9.405 14.470 9.870 14.565 ;
        RECT 9.420 14.460 9.870 14.470 ;
        RECT 6.935 14.205 7.195 14.310 ;
        RECT 5.160 14.035 7.195 14.205 ;
        RECT 5.160 13.960 5.590 14.035 ;
        RECT 2.725 12.730 3.145 12.740 ;
        RECT 4.215 12.730 4.395 13.660 ;
        RECT 1.850 12.550 4.395 12.730 ;
        RECT 2.725 12.280 3.145 12.550 ;
        RECT 5.320 12.150 5.590 13.960 ;
        RECT 6.935 13.950 7.195 14.035 ;
        RECT 7.795 13.940 8.055 14.300 ;
        RECT 10.335 14.275 10.505 15.585 ;
        RECT 11.645 14.275 11.815 15.585 ;
        RECT 12.960 14.275 13.130 15.585 ;
        RECT 14.275 14.275 14.445 15.585 ;
        RECT 15.590 14.275 15.760 15.585 ;
        RECT 16.905 14.275 17.075 15.585 ;
        RECT 18.220 14.275 18.390 15.585 ;
        RECT 5.855 13.845 6.115 13.890 ;
        RECT 5.855 13.800 6.215 13.845 ;
        RECT 7.840 13.800 8.010 13.940 ;
        RECT 10.285 13.915 10.545 14.275 ;
        RECT 11.595 13.915 11.855 14.275 ;
        RECT 12.910 13.915 13.170 14.275 ;
        RECT 14.225 13.915 14.485 14.275 ;
        RECT 15.540 13.915 15.800 14.275 ;
        RECT 16.855 13.915 17.115 14.275 ;
        RECT 18.170 13.915 18.430 14.275 ;
        RECT 5.855 13.630 8.010 13.800 ;
        RECT 5.855 13.585 6.215 13.630 ;
        RECT 5.855 13.530 6.115 13.585 ;
        RECT 7.185 13.110 7.445 13.210 ;
        RECT 9.455 13.110 9.730 13.160 ;
        RECT 7.185 12.940 9.730 13.110 ;
        RECT 7.185 12.850 7.445 12.940 ;
        RECT 9.455 12.900 9.730 12.940 ;
        RECT 5.320 11.890 19.840 12.150 ;
        RECT 7.620 3.690 10.450 11.470 ;
        RECT 14.340 7.200 17.170 10.830 ;
        RECT 19.580 7.590 19.840 11.890 ;
        RECT 20.500 9.040 20.760 23.040 ;
        RECT 24.400 22.990 32.280 23.040 ;
        RECT 29.300 21.450 31.270 21.820 ;
        RECT 27.830 21.070 28.090 21.410 ;
        RECT 33.040 21.070 33.300 24.600 ;
        RECT 34.065 24.325 36.870 26.150 ;
        RECT 34.060 23.300 41.940 23.350 ;
        RECT 34.060 23.040 45.980 23.300 ;
        RECT 34.060 22.990 41.940 23.040 ;
        RECT 35.300 21.450 37.270 21.820 ;
        RECT 38.470 21.070 38.730 21.410 ;
        RECT 27.830 20.810 38.730 21.070 ;
        RECT 27.830 20.470 28.090 20.810 ;
        RECT 33.040 20.800 33.300 20.810 ;
        RECT 28.345 20.130 38.225 20.490 ;
        RECT 38.470 20.470 38.730 20.810 ;
        RECT 31.770 19.645 34.580 20.130 ;
        RECT 22.010 16.620 22.350 19.340 ;
        RECT 25.130 18.590 29.895 18.970 ;
        RECT 22.010 14.570 22.340 16.620 ;
        RECT 22.010 14.220 22.350 14.570 ;
        RECT 22.520 11.520 23.240 17.830 ;
        RECT 23.720 12.660 24.440 16.620 ;
        RECT 31.780 14.570 32.500 19.645 ;
        RECT 32.640 14.220 32.980 19.340 ;
        RECT 33.370 13.130 33.710 16.970 ;
        RECT 33.860 14.550 34.580 19.645 ;
        RECT 24.180 11.940 24.440 12.660 ;
        RECT 41.910 12.330 42.630 16.600 ;
        RECT 41.910 12.280 42.580 12.330 ;
        RECT 27.330 11.940 27.590 11.950 ;
        RECT 41.910 11.940 42.170 12.280 ;
        RECT 24.180 11.680 27.590 11.940 ;
        RECT 27.330 11.520 27.590 11.680 ;
        RECT 38.920 11.680 42.170 11.940 ;
        RECT 38.920 11.520 39.180 11.680 ;
        RECT 43.110 11.520 43.830 17.840 ;
        RECT 44.010 13.130 44.340 16.980 ;
        RECT 21.480 11.160 25.360 11.520 ;
        RECT 27.330 11.160 32.210 11.520 ;
        RECT 34.300 11.160 39.180 11.520 ;
        RECT 40.980 11.160 44.860 11.520 ;
        RECT 27.330 9.040 32.210 9.090 ;
        RECT 20.500 8.780 32.210 9.040 ;
        RECT 27.330 8.730 32.210 8.780 ;
        RECT 32.410 7.790 32.670 11.160 ;
        RECT 33.840 7.790 34.100 11.160 ;
        RECT 34.300 9.040 39.180 9.090 ;
        RECT 45.590 9.040 45.850 23.040 ;
        RECT 34.300 8.780 45.850 9.040 ;
        RECT 34.300 8.730 39.180 8.780 ;
        RECT 34.770 7.590 35.030 8.730 ;
        RECT 19.580 7.330 35.030 7.590 ;
        RECT 20.540 6.800 45.800 7.180 ;
        RECT 7.620 2.200 8.340 3.690 ;
        RECT 7.620 1.380 13.490 2.200 ;
      LAYER via2 ;
        RECT 5.180 50.840 5.550 52.070 ;
        RECT 7.060 50.940 7.430 52.170 ;
        RECT 18.520 46.640 20.530 47.000 ;
        RECT 22.100 45.690 24.110 46.050 ;
        RECT 20.545 43.340 45.805 43.620 ;
        RECT 12.630 42.330 17.510 42.610 ;
        RECT 6.970 26.650 17.840 26.930 ;
        RECT 15.960 24.390 18.010 25.330 ;
        RECT 29.345 28.690 31.225 28.970 ;
        RECT 35.345 28.690 37.225 28.970 ;
        RECT 6.200 17.355 18.825 17.635 ;
        RECT 14.420 7.330 17.070 7.610 ;
        RECT 29.345 21.500 31.225 21.780 ;
        RECT 34.065 24.375 36.870 26.100 ;
        RECT 35.345 21.500 37.225 21.780 ;
        RECT 25.130 18.640 29.895 18.920 ;
        RECT 20.540 6.850 45.800 7.130 ;
        RECT 7.620 1.430 13.490 2.150 ;
      LAYER met3 ;
        RECT 5.130 50.815 5.600 52.095 ;
        RECT 7.010 50.915 7.480 52.195 ;
        RECT 18.470 46.615 20.580 47.025 ;
        RECT 22.050 45.665 24.160 46.075 ;
        RECT 1.320 45.365 1.780 45.370 ;
        RECT 1.320 45.360 45.985 45.365 ;
        RECT 1.320 43.320 50.495 45.360 ;
        RECT 1.630 43.315 50.495 43.320 ;
        RECT 12.630 42.635 17.510 43.315 ;
        RECT 12.580 42.305 17.560 42.635 ;
        RECT 3.855 33.560 37.225 33.565 ;
        RECT 1.000 31.565 37.225 33.560 ;
        RECT 1.000 26.955 5.220 31.565 ;
        RECT 29.345 28.995 31.225 31.565 ;
        RECT 35.345 28.995 37.225 31.565 ;
        RECT 29.295 28.665 31.275 28.995 ;
        RECT 35.295 28.665 37.275 28.995 ;
        RECT 1.000 26.290 17.890 26.955 ;
        RECT 29.345 26.290 31.225 28.665 ;
        RECT 35.345 26.550 37.225 28.665 ;
        RECT 35.345 26.290 37.220 26.550 ;
        RECT 1.000 24.200 37.220 26.290 ;
        RECT 1.000 24.190 37.225 24.200 ;
        RECT 1.000 18.910 5.220 24.190 ;
        RECT 29.345 21.805 31.225 24.190 ;
        RECT 35.345 21.805 37.225 24.190 ;
        RECT 29.295 21.475 31.275 21.805 ;
        RECT 35.295 21.475 37.275 21.805 ;
        RECT 29.345 18.945 31.225 21.475 ;
        RECT 25.080 18.910 31.225 18.945 ;
        RECT 35.345 19.100 37.225 21.475 ;
        RECT 35.345 18.910 37.220 19.100 ;
        RECT 1.000 16.910 37.220 18.910 ;
        RECT 14.340 7.155 17.170 7.640 ;
        RECT 43.985 7.155 50.495 43.315 ;
        RECT 1.410 7.105 2.540 7.110 ;
        RECT 6.255 7.105 50.495 7.155 ;
        RECT 1.410 5.110 50.495 7.105 ;
        RECT 1.470 5.105 50.495 5.110 ;
        RECT 43.985 5.000 50.495 5.105 ;
        RECT 7.570 1.405 13.540 2.175 ;
      LAYER via3 ;
        RECT 5.180 50.840 5.550 52.070 ;
        RECT 7.060 50.940 7.430 52.170 ;
        RECT 18.520 46.640 20.530 47.000 ;
        RECT 22.100 45.690 24.110 46.050 ;
        RECT 1.100 17.010 2.400 33.460 ;
        RECT 49.095 5.100 50.395 45.260 ;
        RECT 7.620 1.430 13.490 2.150 ;
      LAYER met4 ;
        RECT 147.475 224.760 147.510 225.760 ;
        RECT 147.810 224.765 147.840 225.760 ;
        RECT 147.810 224.760 147.845 224.765 ;
        RECT 88.630 224.170 88.930 224.760 ;
        RECT 88.590 223.295 88.975 224.170 ;
        RECT 5.180 222.925 88.975 223.295 ;
        RECT 5.180 52.075 5.550 222.925 ;
        RECT 147.475 222.585 147.845 224.760 ;
        RECT 7.060 222.215 147.845 222.585 ;
        RECT 7.060 52.175 7.430 222.215 ;
        RECT 5.175 50.835 5.555 52.075 ;
        RECT 7.055 50.935 7.435 52.175 ;
        RECT 18.515 47.000 20.535 47.005 ;
        RECT 18.515 46.640 48.630 47.000 ;
        RECT 18.515 46.635 20.535 46.640 ;
        RECT 22.095 46.050 24.115 46.055 ;
        RECT 22.095 45.690 47.260 46.050 ;
        RECT 22.095 45.685 24.115 45.690 ;
        RECT 46.900 3.200 47.260 45.690 ;
        RECT 48.270 4.470 48.630 46.640 ;
        RECT 48.270 4.110 157.040 4.470 ;
        RECT 46.900 2.840 134.950 3.200 ;
        RECT 7.615 2.150 13.495 2.155 ;
        RECT 7.615 1.430 113.060 2.150 ;
        RECT 7.615 1.425 13.495 1.430 ;
        RECT 112.340 1.000 113.060 1.430 ;
        RECT 134.590 1.000 134.950 2.840 ;
        RECT 156.680 1.000 157.040 4.110 ;
        RECT 112.340 0.680 112.400 1.000 ;
        RECT 113.000 0.680 113.060 1.000 ;
  END
END tt_um_vaf_555_timer
END LIBRARY

