magic
tech sky130A
magscale 1 2
timestamp 1711728332
<< pwell >>
rect -106 -170 104 102
<< nmos >>
rect -15 -131 15 69
<< ndiff >>
rect -73 57 -15 69
rect -73 -119 -61 57
rect -27 -119 -15 57
rect -73 -131 -15 -119
rect 15 57 73 69
rect 15 -120 27 57
rect 61 -120 73 57
rect 15 -131 73 -120
<< ndiffc >>
rect -61 -119 -27 57
rect 27 -120 61 57
<< poly >>
rect -15 69 15 95
rect -15 -157 15 -131
<< locali >>
rect -61 57 -27 73
rect 27 57 61 73
rect -61 -135 -27 -119
rect 25 -120 27 57
rect 61 -120 63 57
rect 25 -136 63 -120
<< viali >>
rect -61 -119 -27 57
rect 27 -120 61 57
<< metal1 >>
rect -67 57 -21 69
rect -67 -119 -61 57
rect -27 -119 -21 57
rect -67 -131 -21 -119
rect 21 57 67 69
rect 21 -120 27 57
rect 61 -120 67 57
rect 21 -132 67 -120
<< properties >>
string FIXED_BBOX -158 -226 158 226
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
