magic
tech sky130A
magscale 1 2
timestamp 1711855675
<< error_p >>
rect -287 1072 -225 1078
rect -159 1072 -97 1078
rect -31 1072 31 1078
rect 97 1072 159 1078
rect 225 1072 287 1078
rect -287 1038 -275 1072
rect -159 1038 -147 1072
rect -31 1038 -19 1072
rect 97 1038 109 1072
rect 225 1038 237 1072
rect -287 1032 -225 1038
rect -159 1032 -97 1038
rect -31 1032 31 1038
rect 97 1032 159 1038
rect 225 1032 287 1038
rect -287 -1038 -225 -1032
rect -159 -1038 -97 -1032
rect -31 -1038 31 -1032
rect 97 -1038 159 -1032
rect 225 -1038 287 -1032
rect -287 -1072 -275 -1038
rect -159 -1072 -147 -1038
rect -31 -1072 -19 -1038
rect 97 -1072 109 -1038
rect 225 -1072 237 -1038
rect -287 -1078 -225 -1072
rect -159 -1078 -97 -1072
rect -31 -1078 31 -1072
rect 97 -1078 159 -1072
rect 225 -1078 287 -1072
<< pwell >>
rect -487 -1210 487 1210
<< nmoslvt >>
rect -291 -1000 -221 1000
rect -163 -1000 -93 1000
rect -35 -1000 35 1000
rect 93 -1000 163 1000
rect 221 -1000 291 1000
<< ndiff >>
rect -349 988 -291 1000
rect -349 -988 -337 988
rect -303 -988 -291 988
rect -349 -1000 -291 -988
rect -221 988 -163 1000
rect -221 -988 -209 988
rect -175 -988 -163 988
rect -221 -1000 -163 -988
rect -93 988 -35 1000
rect -93 -988 -81 988
rect -47 -988 -35 988
rect -93 -1000 -35 -988
rect 35 988 93 1000
rect 35 -988 47 988
rect 81 -988 93 988
rect 35 -1000 93 -988
rect 163 988 221 1000
rect 163 -988 175 988
rect 209 -988 221 988
rect 163 -1000 221 -988
rect 291 988 349 1000
rect 291 -988 303 988
rect 337 -988 349 988
rect 291 -1000 349 -988
<< ndiffc >>
rect -337 -988 -303 988
rect -209 -988 -175 988
rect -81 -988 -47 988
rect 47 -988 81 988
rect 175 -988 209 988
rect 303 -988 337 988
<< psubdiff >>
rect -451 1140 -355 1174
rect 355 1140 451 1174
rect -451 1078 -417 1140
rect 417 1078 451 1140
rect -451 -1140 -417 -1078
rect 417 -1140 451 -1078
rect -451 -1174 -355 -1140
rect 355 -1174 451 -1140
<< psubdiffcont >>
rect -355 1140 355 1174
rect -451 -1078 -417 1078
rect 417 -1078 451 1078
rect -355 -1174 355 -1140
<< poly >>
rect -291 1072 -221 1088
rect -291 1038 -275 1072
rect -237 1038 -221 1072
rect -291 1000 -221 1038
rect -163 1072 -93 1088
rect -163 1038 -147 1072
rect -109 1038 -93 1072
rect -163 1000 -93 1038
rect -35 1072 35 1088
rect -35 1038 -19 1072
rect 19 1038 35 1072
rect -35 1000 35 1038
rect 93 1072 163 1088
rect 93 1038 109 1072
rect 147 1038 163 1072
rect 93 1000 163 1038
rect 221 1072 291 1088
rect 221 1038 237 1072
rect 275 1038 291 1072
rect 221 1000 291 1038
rect -291 -1038 -221 -1000
rect -291 -1072 -275 -1038
rect -237 -1072 -221 -1038
rect -291 -1088 -221 -1072
rect -163 -1038 -93 -1000
rect -163 -1072 -147 -1038
rect -109 -1072 -93 -1038
rect -163 -1088 -93 -1072
rect -35 -1038 35 -1000
rect -35 -1072 -19 -1038
rect 19 -1072 35 -1038
rect -35 -1088 35 -1072
rect 93 -1038 163 -1000
rect 93 -1072 109 -1038
rect 147 -1072 163 -1038
rect 93 -1088 163 -1072
rect 221 -1038 291 -1000
rect 221 -1072 237 -1038
rect 275 -1072 291 -1038
rect 221 -1088 291 -1072
<< polycont >>
rect -275 1038 -237 1072
rect -147 1038 -109 1072
rect -19 1038 19 1072
rect 109 1038 147 1072
rect 237 1038 275 1072
rect -275 -1072 -237 -1038
rect -147 -1072 -109 -1038
rect -19 -1072 19 -1038
rect 109 -1072 147 -1038
rect 237 -1072 275 -1038
<< locali >>
rect -451 1140 -355 1174
rect 355 1140 451 1174
rect -451 1078 -417 1140
rect 417 1078 451 1140
rect -291 1038 -275 1072
rect -237 1038 -221 1072
rect -163 1038 -147 1072
rect -109 1038 -93 1072
rect -35 1038 -19 1072
rect 19 1038 35 1072
rect 93 1038 109 1072
rect 147 1038 163 1072
rect 221 1038 237 1072
rect 275 1038 291 1072
rect -337 988 -303 1004
rect -337 -1004 -303 -988
rect -209 988 -175 1004
rect -209 -1004 -175 -988
rect -81 988 -47 1004
rect -81 -1004 -47 -988
rect 47 988 81 1004
rect 47 -1004 81 -988
rect 175 988 209 1004
rect 175 -1004 209 -988
rect 303 988 337 1004
rect 303 -1004 337 -988
rect -291 -1072 -275 -1038
rect -237 -1072 -221 -1038
rect -163 -1072 -147 -1038
rect -109 -1072 -93 -1038
rect -35 -1072 -19 -1038
rect 19 -1072 35 -1038
rect 93 -1072 109 -1038
rect 147 -1072 163 -1038
rect 221 -1072 237 -1038
rect 275 -1072 291 -1038
rect -451 -1140 -417 -1078
rect 417 -1140 451 -1078
rect -451 -1174 -355 -1140
rect 355 -1174 451 -1140
<< viali >>
rect -275 1038 -237 1072
rect -147 1038 -109 1072
rect -19 1038 19 1072
rect 109 1038 147 1072
rect 237 1038 275 1072
rect -337 -988 -303 988
rect -209 -988 -175 988
rect -81 -988 -47 988
rect 47 -988 81 988
rect 175 -988 209 988
rect 303 -988 337 988
rect -275 -1072 -237 -1038
rect -147 -1072 -109 -1038
rect -19 -1072 19 -1038
rect 109 -1072 147 -1038
rect 237 -1072 275 -1038
<< metal1 >>
rect -287 1072 -225 1078
rect -287 1038 -275 1072
rect -237 1038 -225 1072
rect -287 1032 -225 1038
rect -159 1072 -97 1078
rect -159 1038 -147 1072
rect -109 1038 -97 1072
rect -159 1032 -97 1038
rect -31 1072 31 1078
rect -31 1038 -19 1072
rect 19 1038 31 1072
rect -31 1032 31 1038
rect 97 1072 159 1078
rect 97 1038 109 1072
rect 147 1038 159 1072
rect 97 1032 159 1038
rect 225 1072 287 1078
rect 225 1038 237 1072
rect 275 1038 287 1072
rect 225 1032 287 1038
rect -343 988 -297 1000
rect -343 -988 -337 988
rect -303 -988 -297 988
rect -343 -1000 -297 -988
rect -215 988 -169 1000
rect -215 -988 -209 988
rect -175 -988 -169 988
rect -215 -1000 -169 -988
rect -87 988 -41 1000
rect -87 -988 -81 988
rect -47 -988 -41 988
rect -87 -1000 -41 -988
rect 41 988 87 1000
rect 41 -988 47 988
rect 81 -988 87 988
rect 41 -1000 87 -988
rect 169 988 215 1000
rect 169 -988 175 988
rect 209 -988 215 988
rect 169 -1000 215 -988
rect 297 988 343 1000
rect 297 -988 303 988
rect 337 -988 343 988
rect 297 -1000 343 -988
rect -287 -1038 -225 -1032
rect -287 -1072 -275 -1038
rect -237 -1072 -225 -1038
rect -287 -1078 -225 -1072
rect -159 -1038 -97 -1032
rect -159 -1072 -147 -1038
rect -109 -1072 -97 -1038
rect -159 -1078 -97 -1072
rect -31 -1038 31 -1032
rect -31 -1072 -19 -1038
rect 19 -1072 31 -1038
rect -31 -1078 31 -1072
rect 97 -1038 159 -1032
rect 97 -1072 109 -1038
rect 147 -1072 159 -1038
rect 97 -1078 159 -1072
rect 225 -1038 287 -1032
rect 225 -1072 237 -1038
rect 275 -1072 287 -1038
rect 225 -1078 287 -1072
<< properties >>
string FIXED_BBOX -434 -1157 434 1157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 10 l 0.35 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
