magic
tech sky130A
magscale 1 2
timestamp 1711681003
<< error_p >>
rect -479 197 -417 203
rect -351 197 -289 203
rect -223 197 -161 203
rect -95 197 -33 203
rect 33 197 95 203
rect 161 197 223 203
rect 289 197 351 203
rect 417 197 479 203
rect -479 163 -467 197
rect -351 163 -339 197
rect -223 163 -211 197
rect -95 163 -83 197
rect 33 163 45 197
rect 161 163 173 197
rect 289 163 301 197
rect 417 163 429 197
rect -479 157 -417 163
rect -351 157 -289 163
rect -223 157 -161 163
rect -95 157 -33 163
rect 33 157 95 163
rect 161 157 223 163
rect 289 157 351 163
rect 417 157 479 163
rect -479 -163 -417 -157
rect -351 -163 -289 -157
rect -223 -163 -161 -157
rect -95 -163 -33 -157
rect 33 -163 95 -157
rect 161 -163 223 -157
rect 289 -163 351 -157
rect 417 -163 479 -157
rect -479 -197 -467 -163
rect -351 -197 -339 -163
rect -223 -197 -211 -163
rect -95 -197 -83 -163
rect 33 -197 45 -163
rect 161 -197 173 -163
rect 289 -197 301 -163
rect 417 -197 429 -163
rect -479 -203 -417 -197
rect -351 -203 -289 -197
rect -223 -203 -161 -197
rect -95 -203 -33 -197
rect 33 -203 95 -197
rect 161 -203 223 -197
rect 289 -203 351 -197
rect 417 -203 479 -197
<< pwell >>
rect -679 -335 679 335
<< nmoslvt >>
rect -483 -125 -413 125
rect -355 -125 -285 125
rect -227 -125 -157 125
rect -99 -125 -29 125
rect 29 -125 99 125
rect 157 -125 227 125
rect 285 -125 355 125
rect 413 -125 483 125
<< ndiff >>
rect -541 113 -483 125
rect -541 -113 -529 113
rect -495 -113 -483 113
rect -541 -125 -483 -113
rect -413 113 -355 125
rect -413 -113 -401 113
rect -367 -113 -355 113
rect -413 -125 -355 -113
rect -285 113 -227 125
rect -285 -113 -273 113
rect -239 -113 -227 113
rect -285 -125 -227 -113
rect -157 113 -99 125
rect -157 -113 -145 113
rect -111 -113 -99 113
rect -157 -125 -99 -113
rect -29 113 29 125
rect -29 -113 -17 113
rect 17 -113 29 113
rect -29 -125 29 -113
rect 99 113 157 125
rect 99 -113 111 113
rect 145 -113 157 113
rect 99 -125 157 -113
rect 227 113 285 125
rect 227 -113 239 113
rect 273 -113 285 113
rect 227 -125 285 -113
rect 355 113 413 125
rect 355 -113 367 113
rect 401 -113 413 113
rect 355 -125 413 -113
rect 483 113 541 125
rect 483 -113 495 113
rect 529 -113 541 113
rect 483 -125 541 -113
<< ndiffc >>
rect -529 -113 -495 113
rect -401 -113 -367 113
rect -273 -113 -239 113
rect -145 -113 -111 113
rect -17 -113 17 113
rect 111 -113 145 113
rect 239 -113 273 113
rect 367 -113 401 113
rect 495 -113 529 113
<< psubdiff >>
rect -643 265 -547 299
rect 547 265 643 299
rect -643 203 -609 265
rect 609 203 643 265
rect -643 -265 -609 -203
rect 609 -265 643 -203
rect -643 -299 -547 -265
rect 547 -299 643 -265
<< psubdiffcont >>
rect -547 265 547 299
rect -643 -203 -609 203
rect 609 -203 643 203
rect -547 -299 547 -265
<< poly >>
rect -483 197 -413 213
rect -483 163 -467 197
rect -429 163 -413 197
rect -483 125 -413 163
rect -355 197 -285 213
rect -355 163 -339 197
rect -301 163 -285 197
rect -355 125 -285 163
rect -227 197 -157 213
rect -227 163 -211 197
rect -173 163 -157 197
rect -227 125 -157 163
rect -99 197 -29 213
rect -99 163 -83 197
rect -45 163 -29 197
rect -99 125 -29 163
rect 29 197 99 213
rect 29 163 45 197
rect 83 163 99 197
rect 29 125 99 163
rect 157 197 227 213
rect 157 163 173 197
rect 211 163 227 197
rect 157 125 227 163
rect 285 197 355 213
rect 285 163 301 197
rect 339 163 355 197
rect 285 125 355 163
rect 413 197 483 213
rect 413 163 429 197
rect 467 163 483 197
rect 413 125 483 163
rect -483 -163 -413 -125
rect -483 -197 -467 -163
rect -429 -197 -413 -163
rect -483 -213 -413 -197
rect -355 -163 -285 -125
rect -355 -197 -339 -163
rect -301 -197 -285 -163
rect -355 -213 -285 -197
rect -227 -163 -157 -125
rect -227 -197 -211 -163
rect -173 -197 -157 -163
rect -227 -213 -157 -197
rect -99 -163 -29 -125
rect -99 -197 -83 -163
rect -45 -197 -29 -163
rect -99 -213 -29 -197
rect 29 -163 99 -125
rect 29 -197 45 -163
rect 83 -197 99 -163
rect 29 -213 99 -197
rect 157 -163 227 -125
rect 157 -197 173 -163
rect 211 -197 227 -163
rect 157 -213 227 -197
rect 285 -163 355 -125
rect 285 -197 301 -163
rect 339 -197 355 -163
rect 285 -213 355 -197
rect 413 -163 483 -125
rect 413 -197 429 -163
rect 467 -197 483 -163
rect 413 -213 483 -197
<< polycont >>
rect -467 163 -429 197
rect -339 163 -301 197
rect -211 163 -173 197
rect -83 163 -45 197
rect 45 163 83 197
rect 173 163 211 197
rect 301 163 339 197
rect 429 163 467 197
rect -467 -197 -429 -163
rect -339 -197 -301 -163
rect -211 -197 -173 -163
rect -83 -197 -45 -163
rect 45 -197 83 -163
rect 173 -197 211 -163
rect 301 -197 339 -163
rect 429 -197 467 -163
<< locali >>
rect -643 265 -547 299
rect 547 265 643 299
rect -643 203 -609 265
rect 609 203 643 265
rect -483 163 -467 197
rect -429 163 -413 197
rect -355 163 -339 197
rect -301 163 -285 197
rect -227 163 -211 197
rect -173 163 -157 197
rect -99 163 -83 197
rect -45 163 -29 197
rect 29 163 45 197
rect 83 163 99 197
rect 157 163 173 197
rect 211 163 227 197
rect 285 163 301 197
rect 339 163 355 197
rect 413 163 429 197
rect 467 163 483 197
rect -529 113 -495 129
rect -529 -129 -495 -113
rect -401 113 -367 129
rect -401 -129 -367 -113
rect -273 113 -239 129
rect -273 -129 -239 -113
rect -145 113 -111 129
rect -145 -129 -111 -113
rect -17 113 17 129
rect -17 -129 17 -113
rect 111 113 145 129
rect 111 -129 145 -113
rect 239 113 273 129
rect 239 -129 273 -113
rect 367 113 401 129
rect 367 -129 401 -113
rect 495 113 529 129
rect 495 -129 529 -113
rect -483 -197 -467 -163
rect -429 -197 -413 -163
rect -355 -197 -339 -163
rect -301 -197 -285 -163
rect -227 -197 -211 -163
rect -173 -197 -157 -163
rect -99 -197 -83 -163
rect -45 -197 -29 -163
rect 29 -197 45 -163
rect 83 -197 99 -163
rect 157 -197 173 -163
rect 211 -197 227 -163
rect 285 -197 301 -163
rect 339 -197 355 -163
rect 413 -197 429 -163
rect 467 -197 483 -163
rect -643 -265 -609 -203
rect 609 -265 643 -203
rect -643 -299 -547 -265
rect 547 -299 643 -265
<< viali >>
rect -467 163 -429 197
rect -339 163 -301 197
rect -211 163 -173 197
rect -83 163 -45 197
rect 45 163 83 197
rect 173 163 211 197
rect 301 163 339 197
rect 429 163 467 197
rect -529 -113 -495 113
rect -401 -113 -367 113
rect -273 -113 -239 113
rect -145 -113 -111 113
rect -17 -113 17 113
rect 111 -113 145 113
rect 239 -113 273 113
rect 367 -113 401 113
rect 495 -113 529 113
rect -467 -197 -429 -163
rect -339 -197 -301 -163
rect -211 -197 -173 -163
rect -83 -197 -45 -163
rect 45 -197 83 -163
rect 173 -197 211 -163
rect 301 -197 339 -163
rect 429 -197 467 -163
<< metal1 >>
rect -479 197 -417 203
rect -479 163 -467 197
rect -429 163 -417 197
rect -479 157 -417 163
rect -351 197 -289 203
rect -351 163 -339 197
rect -301 163 -289 197
rect -351 157 -289 163
rect -223 197 -161 203
rect -223 163 -211 197
rect -173 163 -161 197
rect -223 157 -161 163
rect -95 197 -33 203
rect -95 163 -83 197
rect -45 163 -33 197
rect -95 157 -33 163
rect 33 197 95 203
rect 33 163 45 197
rect 83 163 95 197
rect 33 157 95 163
rect 161 197 223 203
rect 161 163 173 197
rect 211 163 223 197
rect 161 157 223 163
rect 289 197 351 203
rect 289 163 301 197
rect 339 163 351 197
rect 289 157 351 163
rect 417 197 479 203
rect 417 163 429 197
rect 467 163 479 197
rect 417 157 479 163
rect -535 113 -489 125
rect -535 -113 -529 113
rect -495 -113 -489 113
rect -535 -125 -489 -113
rect -407 113 -361 125
rect -407 -113 -401 113
rect -367 -113 -361 113
rect -407 -125 -361 -113
rect -279 113 -233 125
rect -279 -113 -273 113
rect -239 -113 -233 113
rect -279 -125 -233 -113
rect -151 113 -105 125
rect -151 -113 -145 113
rect -111 -113 -105 113
rect -151 -125 -105 -113
rect -23 113 23 125
rect -23 -113 -17 113
rect 17 -113 23 113
rect -23 -125 23 -113
rect 105 113 151 125
rect 105 -113 111 113
rect 145 -113 151 113
rect 105 -125 151 -113
rect 233 113 279 125
rect 233 -113 239 113
rect 273 -113 279 113
rect 233 -125 279 -113
rect 361 113 407 125
rect 361 -113 367 113
rect 401 -113 407 113
rect 361 -125 407 -113
rect 489 113 535 125
rect 489 -113 495 113
rect 529 -113 535 113
rect 489 -125 535 -113
rect -479 -163 -417 -157
rect -479 -197 -467 -163
rect -429 -197 -417 -163
rect -479 -203 -417 -197
rect -351 -163 -289 -157
rect -351 -197 -339 -163
rect -301 -197 -289 -163
rect -351 -203 -289 -197
rect -223 -163 -161 -157
rect -223 -197 -211 -163
rect -173 -197 -161 -163
rect -223 -203 -161 -197
rect -95 -163 -33 -157
rect -95 -197 -83 -163
rect -45 -197 -33 -163
rect -95 -203 -33 -197
rect 33 -163 95 -157
rect 33 -197 45 -163
rect 83 -197 95 -163
rect 33 -203 95 -197
rect 161 -163 223 -157
rect 161 -197 173 -163
rect 211 -197 223 -163
rect 161 -203 223 -197
rect 289 -163 351 -157
rect 289 -197 301 -163
rect 339 -197 351 -163
rect 289 -203 351 -197
rect 417 -163 479 -157
rect 417 -197 429 -163
rect 467 -197 479 -163
rect 417 -203 479 -197
<< properties >>
string FIXED_BBOX -626 -282 626 282
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.25 l 0.35 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
