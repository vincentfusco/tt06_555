magic
tech sky130A
magscale 1 2
timestamp 1711908466
<< nwell >>
rect 20680 18281 23158 18315
<< pwell >>
rect 20680 17271 23166 17305
<< psubdiff >>
rect 20680 17271 23166 17305
<< nsubdiff >>
rect 24103 19828 28001 19886
rect 20680 18281 23158 18315
<< locali >>
rect 21942 23276 22918 23410
rect 21852 22844 23008 22938
rect 19999 17305 21315 17306
rect 19999 17272 23156 17305
rect 20679 17190 23156 17272
rect 20679 17156 20810 17190
rect 22966 17156 23156 17190
<< viali >>
rect 20810 20140 22984 20174
rect 20810 17156 22966 17190
rect 20696 16384 20748 17094
<< metal1 >>
rect 21932 23276 21942 23332
rect 22918 23276 22928 23332
rect 22962 23062 23030 23080
rect 20798 21930 21230 22720
rect 22598 22438 23030 23062
rect 20798 20914 21230 21704
rect 22598 21422 23030 22212
rect 22598 20514 23030 21196
rect 23120 21088 23172 23884
rect 23330 23184 23382 23884
rect 23515 23478 23525 23534
rect 28577 23478 28587 23534
rect 23320 23132 23330 23184
rect 23382 23132 23392 23184
rect 23246 22282 23322 22288
rect 23246 22224 23252 22282
rect 23316 22279 23322 22282
rect 23316 22227 23498 22279
rect 23316 22224 23322 22227
rect 23246 22218 23322 22224
rect 23120 21036 23544 21088
rect 25275 20548 25285 20604
rect 25661 20548 25671 20604
rect 26475 20548 26485 20604
rect 26861 20548 26871 20604
rect 22938 20368 23030 20514
rect 23352 20372 23428 20378
rect 23352 20368 23358 20372
rect 22938 20316 23358 20368
rect 22938 20304 23030 20316
rect 23352 20314 23358 20316
rect 23422 20314 23428 20372
rect 23352 20308 23428 20314
rect 20909 20196 22885 20288
rect 20800 20180 20810 20196
rect 20798 20140 20810 20180
rect 22984 20180 22994 20196
rect 22984 20140 22996 20180
rect 20798 20134 22996 20140
rect 26219 19916 26229 20030
rect 20798 19510 21230 19862
rect 22598 19688 22608 19876
rect 23018 19688 23028 19876
rect 23522 19798 26229 19916
rect 26219 19685 26229 19798
rect 26790 19916 26800 20030
rect 26790 19798 28576 19916
rect 26790 19685 26800 19798
rect 23246 19512 23322 19518
rect 23246 19510 23252 19512
rect 20798 19458 23252 19510
rect 19696 18964 19706 19332
rect 19758 19016 19768 19332
rect 20798 19100 21230 19458
rect 23246 19454 23252 19458
rect 23316 19454 23322 19512
rect 23246 19448 23322 19454
rect 19758 18964 21018 19016
rect 21070 18964 21080 19016
rect 19698 18590 21230 18872
rect 22598 18679 23030 19352
rect 25275 19110 25285 19166
rect 25661 19110 25671 19166
rect 26475 19110 26485 19166
rect 26861 19110 26871 19166
rect 22598 18625 23510 18679
rect 22598 18590 23030 18625
rect 19698 17292 19888 18590
rect 24432 18538 24442 18590
rect 25395 18538 25405 18590
rect 23336 18484 23346 18536
rect 23398 18484 23408 18536
rect 20646 18281 20656 18333
rect 23181 18281 23191 18333
rect 21745 17876 21779 17980
rect 21745 17867 21778 17876
rect 22270 17867 22304 17994
rect 21565 17833 21778 17867
rect 21827 17833 22103 17867
rect 22162 17833 22304 17867
rect 22353 17833 23209 17867
rect 23218 17833 23262 17867
rect 20228 17701 20339 17735
rect 20123 17356 20134 17364
rect 20193 17356 20201 17364
rect 20560 17292 23166 17305
rect 19698 17271 23166 17292
rect 19698 17190 23156 17271
rect 19698 17156 20810 17190
rect 22966 17156 23156 17190
rect 19698 17150 22978 17156
rect 19698 17094 20754 17150
rect 19698 16384 20696 17094
rect 20748 16384 20754 17094
rect 20930 17042 20940 17094
rect 21506 17042 21516 17094
rect 20810 16448 20856 17030
rect 22920 17014 22966 17030
rect 23228 17014 23262 17833
rect 23346 17488 23398 18484
rect 23346 17436 23490 17488
rect 22920 16976 23262 17014
rect 22274 16914 22284 16966
rect 22850 16914 22860 16966
rect 20930 16786 20940 16838
rect 21506 16786 21516 16838
rect 22274 16658 22284 16710
rect 22850 16658 22860 16710
rect 20930 16530 20940 16582
rect 21506 16530 21516 16582
rect 22920 16448 22966 16976
rect 22274 16384 22284 16436
rect 22850 16384 22860 16436
rect 19698 16338 20754 16384
rect 19698 16332 28610 16338
rect 19698 16276 22300 16332
rect 22830 16276 28610 16332
rect 19698 16236 28614 16276
rect 19698 16180 23524 16236
rect 28576 16180 28623 16236
rect 19698 15836 28623 16180
<< via1 >>
rect 21942 23276 22918 23332
rect 23525 23478 28577 23534
rect 23330 23132 23382 23184
rect 23252 22224 23316 22282
rect 25285 20548 25661 20604
rect 26485 20548 26861 20604
rect 23358 20314 23422 20372
rect 20810 20174 22984 20196
rect 20810 20140 22984 20174
rect 22608 19688 23018 19876
rect 26229 19685 26790 20030
rect 19706 18964 19758 19332
rect 23252 19454 23316 19512
rect 21018 18964 21070 19016
rect 25285 19110 25661 19166
rect 26485 19110 26861 19166
rect 24442 18538 25395 18590
rect 23346 18484 23398 18536
rect 20656 18281 23181 18333
rect 20940 17042 21506 17094
rect 22284 16914 22850 16966
rect 20940 16786 21506 16838
rect 22284 16658 22850 16710
rect 20940 16530 21506 16582
rect 22284 16384 22850 16436
rect 22300 16276 22830 16332
rect 23524 16180 28576 16236
<< metal2 >>
rect 19706 19332 19758 23886
rect 19706 18954 19758 18964
rect 19786 17356 19850 23889
rect 23525 23534 28577 23544
rect 23525 23468 28577 23478
rect 19879 23388 28588 23440
rect 19879 17992 19931 23388
rect 21942 23332 22918 23342
rect 21942 23266 22918 23276
rect 23330 23184 23382 23194
rect 23330 22928 23382 23132
rect 28536 23126 28588 23388
rect 23128 22876 23382 22928
rect 20810 20196 22984 20206
rect 20810 20130 22984 20140
rect 22608 19876 23018 19886
rect 22608 19678 23018 19688
rect 23128 19216 23180 22876
rect 23246 22282 23322 22288
rect 23246 22224 23252 22282
rect 23316 22224 23322 22282
rect 23246 22218 23322 22224
rect 23258 19518 23310 22218
rect 25285 20604 25661 20614
rect 25285 20538 25661 20548
rect 26485 20604 26861 20614
rect 26485 20538 26861 20548
rect 23352 20372 23428 20378
rect 23352 20314 23358 20372
rect 23422 20314 23428 20372
rect 23352 20308 23428 20314
rect 23364 19984 23416 20308
rect 26229 20030 26790 20040
rect 23364 19932 23492 19984
rect 23364 19782 23416 19932
rect 23364 19730 23490 19782
rect 26229 19675 26790 19685
rect 23246 19512 23322 19518
rect 23246 19454 23252 19512
rect 23316 19454 23322 19512
rect 23246 19448 23322 19454
rect 23128 19164 23398 19216
rect 21018 19016 21070 19026
rect 21070 18964 23290 19016
rect 21018 18954 21070 18964
rect 20656 18337 23181 18347
rect 20656 18271 23181 18281
rect 19879 17938 20014 17992
rect 23238 17989 23290 18964
rect 23346 18536 23398 19164
rect 25276 19166 25670 19174
rect 25276 19110 25285 19166
rect 25661 19110 25670 19166
rect 25276 19100 25670 19110
rect 26476 19166 26870 19174
rect 26476 19110 26485 19166
rect 26861 19110 26870 19166
rect 26476 19100 26870 19110
rect 24442 18594 25395 18604
rect 24442 18528 25395 18538
rect 23346 18474 23398 18484
rect 21356 17776 21390 17989
rect 23052 17980 23290 17989
rect 21621 17946 21937 17980
rect 22147 17946 23290 17980
rect 23052 17937 23290 17946
rect 23238 17936 23290 17937
rect 19786 17320 20122 17356
rect 20480 17240 20534 17769
rect 21300 17702 21390 17776
rect 21310 17390 21362 17442
rect 20480 17188 23384 17240
rect 20940 17094 21506 17104
rect 20940 16838 21506 17042
rect 20940 16582 21506 16786
rect 20940 15832 21506 16530
rect 22284 16966 22850 16976
rect 22284 16710 22850 16914
rect 22284 16436 22850 16658
rect 22284 16332 22850 16384
rect 22284 16276 22300 16332
rect 22830 16276 22850 16332
rect 23332 16328 23384 17188
rect 26370 16328 26422 16618
rect 23332 16276 26422 16328
rect 22284 16250 22850 16276
rect 23524 16236 28576 16246
rect 23524 16170 28576 16180
<< via2 >>
rect 23525 23478 28577 23534
rect 21942 23276 22918 23332
rect 20810 20140 22984 20196
rect 22608 19688 23018 19876
rect 25285 20548 25661 20604
rect 26485 20548 26861 20604
rect 26229 19685 26790 20030
rect 20656 18333 23181 18337
rect 20656 18281 23181 18333
rect 25285 19110 25661 19166
rect 26485 19110 26861 19166
rect 24442 18590 25395 18594
rect 24442 18538 25395 18590
rect 22300 16276 22830 16332
rect 23524 16180 28576 16236
<< metal3 >>
rect 19680 23883 19772 23884
rect 19680 23534 28613 23883
rect 19680 23478 23525 23534
rect 28577 23478 28613 23534
rect 19680 23474 28613 23478
rect 19742 23473 28613 23474
rect 21942 23337 22918 23473
rect 21932 23332 22928 23337
rect 21932 23276 21942 23332
rect 22918 23276 22928 23332
rect 21932 23271 22928 23276
rect 20187 21522 26861 21523
rect 19697 21123 26861 21522
rect 19697 20201 20167 21123
rect 25285 20609 25661 21123
rect 26485 20609 26861 21123
rect 25275 20604 25671 20609
rect 25275 20548 25285 20604
rect 25661 20548 25671 20604
rect 25275 20543 25671 20548
rect 26475 20604 26871 20609
rect 26475 20548 26485 20604
rect 26861 20548 26871 20604
rect 26475 20543 26871 20548
rect 19697 20196 22994 20201
rect 19697 20140 20810 20196
rect 22984 20140 22994 20196
rect 19697 20068 22994 20140
rect 25285 20068 25661 20543
rect 26485 20120 26861 20543
rect 26485 20068 26860 20120
rect 19697 20030 26860 20068
rect 19697 19876 26229 20030
rect 19697 19688 22608 19876
rect 23018 19688 26229 19876
rect 19697 19685 26229 19688
rect 26790 19685 26860 20030
rect 19697 19650 26860 19685
rect 19697 19648 26861 19650
rect 19697 18592 20167 19648
rect 25285 19171 25661 19648
rect 26485 19171 26861 19648
rect 25275 19166 25671 19171
rect 25275 19110 25285 19166
rect 25661 19110 25671 19166
rect 25275 19105 25671 19110
rect 26475 19166 26871 19171
rect 26475 19110 26485 19166
rect 26861 19110 26871 19166
rect 26475 19105 26871 19110
rect 25285 18599 25661 19105
rect 24432 18594 25661 18599
rect 24432 18592 24442 18594
rect 19697 18538 24442 18592
rect 25395 18592 25661 18594
rect 26485 18630 26861 19105
rect 26485 18592 26860 18630
rect 25395 18538 26860 18592
rect 19697 18337 26860 18538
rect 19697 18281 20656 18337
rect 23181 18281 26860 18337
rect 19697 18193 26860 18281
rect 19765 18192 26860 18193
rect 22284 16332 22850 16338
rect 22284 16276 22300 16332
rect 22830 16276 22850 16332
rect 22284 16241 22850 16276
rect 28213 16241 28613 23473
rect 20667 16236 28613 16241
rect 19698 16231 19924 16232
rect 20667 16231 23524 16236
rect 19698 16180 23524 16231
rect 28576 16180 28613 16236
rect 19698 15894 28613 16180
rect 19698 15832 28623 15894
rect 19710 15831 28623 15832
use comp_p  X_COMP_P_BOTTOM
timestamp 1711855675
transform 1 0 26492 0 1 14702
box -3002 1462 2120 5166
use comp_p  X_COMP_P_TOP
timestamp 1711855675
transform 1 0 26493 0 -1 25012
box -3002 1462 2120 5166
use inv  X_INV1
timestamp 1711908466
transform 1 0 20381 0 1 16477
box 978 788 1260 1874
use inv  X_INV2[0]
timestamp 1711908466
transform 1 0 20906 0 1 16477
box 978 788 1260 1874
use inv  X_INV2[1]
timestamp 1711908466
transform 1 0 20643 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[0]
timestamp 1711908466
transform 1 0 21958 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[1]
timestamp 1711908466
transform 1 0 21695 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[2]
timestamp 1711908466
transform 1 0 21432 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[3]
timestamp 1711908466
transform 1 0 21169 0 1 16477
box 978 788 1260 1874
use sr_latch_rb  X_SR_LATCH
timestamp 1711908466
transform 1 0 26627 0 1 16912
box -6666 354 -5267 1440
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_bias
timestamp 1711855675
transform 0 1 22430 -1 0 23164
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_NVJ7JE  XMn_discharge
timestamp 1711855675
transform 0 1 21888 -1 0 16739
box -487 -1210 487 1210
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_bias
timestamp 1711855675
transform 0 1 21897 -1 0 20400
box -296 -1219 296 1219
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_1
timestamp 1711855675
transform 0 1 21914 1 0 21055
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_2
timestamp 1711855675
transform 0 1 21914 1 0 21563
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_3
timestamp 1711855675
transform 0 1 21914 1 0 22071
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_4
timestamp 1711855675
transform 0 1 21914 1 0 22579
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bot
timestamp 1711855675
transform 0 1 21914 -1 0 18731
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_mid
timestamp 1711855675
transform 0 1 21914 -1 0 19239
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_top
timestamp 1711855675
transform 0 1 21914 -1 0 19747
box -307 -1282 307 1282
<< labels >>
flabel metal1 23120 23832 23172 23884 3 FreeSans 960 270 0 0 V_THRESH_I
port 0 e default input
flabel metal2 20940 15832 21506 15888 1 FreeSans 1280 0 0 0 V_DISCH_O
port 4 n default output
flabel metal3 23524 15836 28576 15892 1 FreeSans 960 0 0 0 VSS
port 6 n default bidirectional
flabel metal1 23330 23832 23382 23884 7 FreeSans 960 90 0 0 V_TRIG_B_I
port 1 w default input
flabel metal1 22828 18724 22828 18724 1 FreeSans 640 0 0 0 v0p6
flabel metal1 21034 19270 21034 19270 1 FreeSans 960 0 0 0 v1p2
flabel metal2 21346 17736 21346 17736 1 FreeSans 320 0 0 0 q_sr
flabel metal1 21672 17852 21674 17852 1 FreeSans 320 0 0 0 out_inv1
flabel metal1 23138 16992 23140 16992 1 FreeSans 320 0 0 0 out_inv3
flabel metal1 22814 22574 22814 22574 1 FreeSans 640 0 0 0 bias_n
flabel metal1 21010 22070 21010 22070 1 FreeSans 640 0 0 0 bias_3
flabel metal1 22812 22072 22812 22072 1 FreeSans 640 0 0 0 bias_2
flabel metal1 21014 21056 21014 21056 1 FreeSans 640 0 0 0 bias_1
flabel metal1 22754 20966 22754 20966 1 FreeSans 640 0 0 0 bias_p
flabel metal2 21338 17416 21338 17418 1 FreeSans 320 0 0 0 qb_sr
flabel metal3 19698 19116 19754 21458 3 FreeSans 960 0 0 0 VDD
port 5 e default bidirectional
flabel metal2 19706 23834 19758 23886 3 FreeSans 960 270 0 0 DO_OUT
port 3 e default output
flabel metal2 19792 23822 19848 23888 7 FreeSans 960 90 0 0 DI_RESET_N
port 2 w default input
<< end >>
