** sch_path: /home/vincef/projects/tt06_555/xsch/ip/timers/timer_core/timer_core.sch
.subckt timer_core V_THRESH_I V_TRIG_B_I DO_OUT V_DISCH_O VDD VSS
*.PININFO V_THRESH_I:I V_TRIG_B_I:I DO_OUT:O VDD:B VSS:B V_DISCH_O:O
XR_top v1p2 VDD VSS sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
XR_mid v0p6 v1p2 VSS sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
XR_bot VSS v0p6 VSS sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
* noconn qb_sr
XR_bias_1 bias_1 bias_p VSS sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
XMn_bias bias_n bias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=1
XMp_bias bias_p bias_p VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=10 nf=1 m=1
XMn_discharge V_DISCH_O out_inv3 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.35 W=10 nf=1 m=5
XR_bias_2 bias_2 bias_1 VSS sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
XR_bias_3 bias_3 bias_2 VSS sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
XR_bias_4 bias_n bias_3 VSS sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
X_INV3[3] DO_OUT out_inv3 VDD VSS inv
X_INV3[2] DO_OUT out_inv3 VDD VSS inv
X_INV3[1] DO_OUT out_inv3 VDD VSS inv
X_INV3[0] DO_OUT out_inv3 VDD VSS inv
X_INV2[1] out_inv1 DO_OUT VDD VSS inv
X_INV2[0] out_inv1 DO_OUT VDD VSS inv
X_INV1 q_sr out_inv1 VDD VSS inv
X_SR_LATCH sr_s qb_sr VDD VSS sr_r q_sr sr_latch
X_COMP_P_BOTTOM v0p6 sr_s VDD VSS V_TRIG_B_I bias_p comp_p
X_COMP_P_TOP V_THRESH_I sr_r VDD VSS v1p2 bias_p comp_p
.ends

* expanding   symbol:  ip/logic/inv/inv.sym # of pins=4
** sym_path: /home/vincef/projects/tt06_555/xsch/ip/logic/inv/inv.sym
** sch_path: /home/vincef/projects/tt06_555/xsch/ip/logic/inv/inv.sch
.subckt inv vin vout vdd vss
*.PININFO vin:I vout:O vdd:I vss:I
XMn vout vin vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XMp vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  ip/logic/sr_latch/sr_latch.sym # of pins=6
** sym_path: /home/vincef/projects/tt06_555/xsch/ip/logic/sr_latch/sr_latch.sym
** sch_path: /home/vincef/projects/tt06_555/xsch/ip/logic/sr_latch/sr_latch.sch
.subckt sr_latch IN_S OUT_Q_B vdd vss IN_R OUT_Q
*.PININFO IN_R:I OUT_Q_B:O OUT_Q:O IN_S:I vdd:I vss:I
X_NOR_TOP OUT_Q OUT_Q_B vdd vss IN_S nor
X_NOR_BOTTOM OUT_Q_B OUT_Q vdd vss IN_R nor
.ends


* expanding   symbol:  ip/comparators/comp_p/comp_p.sym # of pins=6
** sym_path: /home/vincef/projects/tt06_555/xsch/ip/comparators/comp_p/comp_p.sym
** sch_path: /home/vincef/projects/tt06_555/xsch/ip/comparators/comp_p/comp_p.sch
.subckt comp_p vinp vout vdd vss vinn vbias_p
*.PININFO vdd:B vss:B vbias_p:I vinn:I vinp:I vout:O
XMp_inn1 latch_left vinn tail vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 m=4
XMp_inp1 latch_right vinp tail vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 m=4
XMn_diode_left1 latch_left latch_left vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XMn_cs_left latch_right latch_left vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=1
XMn_diode_right latch_right latch_right vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XMn_cs_right1 latch_left latch_right vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=1
XMp_tail tail vbias_p vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=10 nf=1 m=1
XMn_out_right vout latch_right vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=1
XMn_out_left out_left latch_left vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=1
XMp_diode_left1 out_left out_left vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 m=1
XMp_out vout out_left vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 m=1
.ends


* expanding   symbol:  ip/logic/nor/nor.sym # of pins=5
** sym_path: /home/vincef/projects/tt06_555/xsch/ip/logic/nor/nor.sym
** sch_path: /home/vincef/projects/tt06_555/xsch/ip/logic/nor/nor.sch
.subckt nor IN_A OUT vdd vss IN_B
*.PININFO IN_A:I OUT:O vss:B vdd:B IN_B:I
XMn_a OUT IN_A vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XMp_a mpcon IN_A vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XMp_b OUT IN_B mpcon vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XMn_b OUT IN_B vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
