magic
tech sky130A
magscale 1 2
timestamp 1711732688
<< nwell >>
rect 978 1218 1260 1437
<< pwell >>
rect 978 788 1260 1218
<< psubdiff >>
rect 1016 794 1040 828
rect 1198 794 1222 828
<< psubdiffcont >>
rect 1040 794 1198 828
<< poly >>
rect 1104 1453 1134 1504
rect 1086 1169 1152 1185
rect 1086 1135 1102 1169
rect 1136 1135 1152 1169
rect 1086 1119 1152 1135
rect 1104 1082 1134 1119
<< polycont >>
rect 1102 1135 1136 1169
<< locali >>
rect 1086 1135 1102 1169
rect 1136 1135 1152 1169
rect 1024 794 1040 828
rect 1198 794 1214 828
<< viali >>
rect 1040 1804 1198 1838
rect 1102 1135 1136 1169
rect 1040 794 1198 828
<< metal1 >>
rect 1028 1838 1210 1844
rect 1028 1804 1040 1838
rect 1198 1804 1210 1838
rect 1028 1798 1210 1804
rect 1058 1562 1092 1798
rect 1140 1548 1218 1754
rect 1102 1390 1136 1504
rect 978 1356 1136 1390
rect 1102 1186 1136 1356
rect 1184 1390 1218 1548
rect 1184 1356 1260 1390
rect 1085 1169 1152 1186
rect 1085 1135 1102 1169
rect 1136 1135 1152 1169
rect 1085 1118 1152 1135
rect 1184 1070 1218 1356
rect 1058 834 1092 1070
rect 1146 878 1218 1070
rect 1028 828 1210 834
rect 1028 794 1040 828
rect 1198 794 1210 828
rect 1028 788 1210 794
use sky130_fd_pr__pfet_01v8_7PK3FC  sky130_fd_pr__pfet_01v8_7PK3FC_0
timestamp 1711732688
transform 1 0 1119 0 1 1614
box -141 -178 141 260
use sky130_fd_pr__nfet_01v8_BXYDM4  XMn
timestamp 1711732688
transform 1 0 1119 0 1 1013
box -106 -216 104 102
<< labels >>
flabel metal1 1040 1804 1198 1838 0 FreeSans 320 0 0 0 vdd
port 3 nsew default bidirectional
flabel metal1 1226 1356 1260 1390 7 FreeSans 320 0 0 0 vout
port 2 w default output
flabel metal1 978 1356 1012 1390 3 FreeSans 320 0 0 0 vin
port 1 e default input
flabel metal1 1040 794 1198 828 0 FreeSans 320 0 0 0 vss
port 4 nsew default bidirectional
<< end >>
