magic
tech sky130A
magscale 1 2
timestamp 1711855675
<< nwell >>
rect -1198 1512 -823 1620
rect -1199 964 -823 1512
<< pwell >>
rect -1200 962 -823 964
rect -1199 540 -823 962
<< nmos >>
rect -1074 628 -1044 828
rect -986 628 -956 828
<< ndiff >>
rect -1132 816 -1074 828
rect -1132 640 -1120 816
rect -1086 640 -1074 816
rect -1132 628 -1074 640
rect -1044 816 -986 828
rect -1044 639 -1032 816
rect -998 639 -986 816
rect -1044 628 -986 639
rect -956 816 -898 828
rect -956 639 -944 816
rect -910 639 -898 816
rect -956 628 -898 639
<< ndiffc >>
rect -1120 640 -1086 816
rect -1032 639 -998 816
rect -944 639 -910 816
<< psubdiff >>
rect -1163 540 -1138 574
rect -892 540 -868 574
<< nsubdiff >>
rect -1154 1550 -1130 1584
rect -892 1550 -868 1584
<< psubdiffcont >>
rect -1138 540 -892 574
<< nsubdiffcont >>
rect -1130 1550 -892 1584
<< poly >>
rect -1074 1019 -1044 1072
rect -1112 1003 -1044 1019
rect -1112 969 -1096 1003
rect -1062 969 -1044 1003
rect -1112 953 -1044 969
rect -1074 828 -1044 953
rect -986 935 -956 1072
rect -1002 919 -936 935
rect -1002 885 -986 919
rect -952 885 -936 919
rect -1002 869 -936 885
rect -986 866 -952 869
rect -986 828 -956 866
rect -1074 602 -1044 628
rect -986 602 -956 628
<< polycont >>
rect -1096 969 -1062 1003
rect -986 885 -952 919
<< locali >>
rect -1146 1550 -1130 1584
rect -892 1550 -876 1584
rect -1032 1460 -998 1550
rect -1112 1003 -1046 1019
rect -1112 969 -1096 1003
rect -1062 969 -1046 1003
rect -1112 953 -1046 969
rect -1002 885 -986 919
rect -952 885 -936 919
rect -982 866 -948 885
rect -1120 816 -1086 832
rect -1120 624 -1086 640
rect -1032 816 -998 832
rect -944 816 -910 832
rect -1032 622 -998 639
rect -946 639 -944 816
rect -910 639 -908 816
rect -946 623 -908 639
rect -1156 540 -1138 574
rect -892 540 -876 574
<< viali >>
rect -1130 1550 -892 1584
rect -1120 1084 -1086 1460
rect -944 1084 -910 1460
rect -1096 969 -1062 1003
rect -986 885 -952 919
rect -1120 640 -1086 816
rect -944 639 -910 816
rect -1138 540 -892 574
<< metal1 >>
rect -1142 1584 -880 1590
rect -1142 1550 -1130 1584
rect -892 1550 -880 1584
rect -1142 1544 -880 1550
rect -1120 1472 -1086 1476
rect -1126 1460 -1080 1472
rect -1126 1084 -1120 1460
rect -1086 1330 -1080 1460
rect -950 1460 -904 1472
rect -950 1330 -944 1460
rect -1086 1214 -944 1330
rect -1086 1084 -1080 1214
rect -1126 1072 -1080 1084
rect -950 1084 -944 1214
rect -910 1098 -904 1460
rect -910 1084 -877 1098
rect -950 1068 -877 1084
rect -1112 1003 -1046 1019
rect -1199 969 -1096 1003
rect -1062 969 -1046 1003
rect -1112 953 -1046 969
rect -1003 919 -935 936
rect -1199 885 -986 919
rect -952 885 -935 919
rect -1003 868 -935 885
rect -907 838 -877 1068
rect -907 832 -823 838
rect -1126 816 -1080 828
rect -1126 640 -1120 816
rect -1086 640 -1080 816
rect -1126 628 -1080 640
rect -950 816 -823 832
rect -950 639 -944 816
rect -910 802 -823 816
rect -910 639 -904 802
rect -1120 580 -1086 628
rect -950 627 -904 639
rect -1150 574 -880 580
rect -1150 540 -1138 574
rect -892 540 -880 574
rect -1150 534 -880 540
use sky130_fd_pr__pfet_01v8_7P3MHC  sky130_fd_pr__pfet_01v8_7P3MHC_1
timestamp 1711855675
transform -1 0 -972 0 1 1236
box -141 -200 138 276
use sky130_fd_pr__pfet_01v8_7P3MHC  sky130_fd_pr__pfet_01v8_7P3MHC_2
timestamp 1711855675
transform -1 0 -1060 0 1 1236
box -141 -200 138 276
<< labels >>
flabel metal1 -1199 885 -1165 919 3 FreeSans 160 0 0 0 IN_B
port 1 e default input
flabel metal1 -1138 540 -892 574 0 FreeSans 320 0 0 0 vss
port 4 nsew default bidirectional
flabel metal1 -1130 1550 -892 1584 0 FreeSans 320 0 0 0 vdd
port 3 nsew default bidirectional
flabel metal1 -1199 969 -1165 1003 3 FreeSans 160 0 0 0 IN_A
port 0 e default input
flabel ndiffc -1014 728 -1014 728 1 FreeSans 80 0 0 0 drain_mna
flabel metal1 -857 803 -823 837 7 FreeSans 160 0 0 0 OUT
port 2 w default output
<< end >>
