* NGSPICE file created from tt_um_vaf_555_timer_flat.ext - technology: sky130A

.subckt tt_um_vaf_555_timer_flat clk ena rst_n ua[3] ua[4] ua[5] ua[6] ua[7] ui_in[1]
+ ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2]
+ uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2]
+ uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2]
+ uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7] ua[2] ui_in[0] uo_out[0] ua[1] ua[0] VGND
+ VPWR
X0 X_TIMER.out_inv3 uo_out[0].t4 VPWR.t9 VPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 X_TIMER.X_COMP_P_BOTTOM.latch_right.t6 X_TIMER.X_COMP_P_BOTTOM.latch_right.t5 VGND.t32 VGND.t31 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X2 X_TIMER.X_COMP_P_TOP.latch_right.t6 ua[0].t0 X_TIMER.X_COMP_P_TOP.tail.t8 VPWR.t12 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X3 X_TIMER.X_COMP_P_TOP.tail.t4 X_TIMER.bias_p VPWR.t38 VPWR.t37 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X4 VPWR.t36 X_TIMER.bias_p X_TIMER.X_COMP_P_BOTTOM.tail.t8 VPWR.t35 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X5 X_TIMER.qb_sr X_TIMER.X_SR_LATCH.IN_S.t2 VGND.t42 VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X6 X_TIMER.out_inv3 uo_out[0].t5 VGND.t4 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X7 X_TIMER.X_SR_LATCH.IN_S.t1 X_TIMER.X_COMP_P_BOTTOM.latch_right.t7 VGND.t30 VGND.t28 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
X8 X_TIMER.X_SR_LATCH.IN_R.t0 X_TIMER.X_COMP_P_TOP.out_left.t3 VPWR.t22 VPWR.t21 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
X9 VGND X_TIMER.v0p6 VGND.t39 sky130_fd_pr__res_xhigh_po_1p41 l=7
X10 X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B ui_in[0].t0 VPWR.t24 VPWR.t23 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X11 X_TIMER.out_inv3 uo_out[0].t6 VGND.t3 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X12 X_TIMER.bias_1 X_TIMER.bias_2 VGND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=7
X13 X_TIMER.X_COMP_P_BOTTOM.tail.t6 ua[1].t0 X_TIMER.X_COMP_P_BOTTOM.latch_left.t6 VPWR.t1 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X14 X_TIMER.out_inv1 X_TIMER.q_sr VPWR.t18 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X15 X_TIMER.X_COMP_P_TOP.latch_right.t5 ua[0].t1 X_TIMER.X_COMP_P_TOP.tail.t6 VPWR.t11 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X16 VPWR.t26 X_TIMER.X_COMP_P_BOTTOM.out_left.t3 X_TIMER.X_SR_LATCH.IN_S.t0 VPWR.t25 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
X17 X_TIMER.out_inv1 X_TIMER.q_sr VGND.t15 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X18 X_TIMER.X_COMP_P_BOTTOM.latch_left.t0 X_TIMER.X_COMP_P_BOTTOM.latch_right.t8 VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
X19 VGND.t13 X_TIMER.X_COMP_P_TOP.latch_left.t7 X_TIMER.X_COMP_P_TOP.out_left.t2 VGND.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
X20 X_TIMER.X_COMP_P_TOP.latch_left.t3 X_TIMER.v1p2 X_TIMER.X_COMP_P_TOP.tail.t1 VPWR.t11 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X21 X_TIMER.bias_p X_TIMER.bias_p VPWR.t34 VPWR.t33 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X22 X_TIMER.X_COMP_P_BOTTOM.tail.t7 ua[1].t1 X_TIMER.X_COMP_P_BOTTOM.latch_left.t5 VPWR.t1 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X23 X_TIMER.X_COMP_P_TOP.latch_left.t2 X_TIMER.v1p2 X_TIMER.X_COMP_P_TOP.tail.t0 VPWR.t12 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X24 X_TIMER.out_inv3 uo_out[0].t7 VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X25 X_TIMER.v1p2 X_TIMER.v0p6 VGND.t39 sky130_fd_pr__res_xhigh_po_1p41 l=7
X26 X_TIMER.X_COMP_P_TOP.latch_left.t1 X_TIMER.v1p2 X_TIMER.X_COMP_P_TOP.tail.t3 VPWR.t11 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X27 X_TIMER.X_SR_LATCH.nand_0.IN_A X_TIMER.X_SR_LATCH.IN_R.t2 VPWR.t14 VPWR.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X28 uo_out[0].t1 X_TIMER.out_inv1 VPWR.t32 VPWR.t31 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X29 X_TIMER.out_inv3 uo_out[0].t8 VPWR.t5 VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X30 X_TIMER.out_inv3 uo_out[0].t9 VGND.t2 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X31 X_TIMER.X_COMP_P_BOTTOM.tail.t3 X_TIMER.v0p6 X_TIMER.X_COMP_P_BOTTOM.latch_right.t3 VPWR.t1 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X32 uo_out[0].t2 X_TIMER.out_inv1 VPWR.t30 VPWR.t29 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X33 VGND.t44 X_TIMER.bias_n X_TIMER.bias_n VGND.t43 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
X34 X_TIMER.q_sr X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B a_1723_2994# VPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X35 X_TIMER.X_COMP_P_BOTTOM.tail.t2 X_TIMER.v0p6 X_TIMER.X_COMP_P_BOTTOM.latch_right.t2 VPWR.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X36 X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B ui_in[0].t1 X_TIMER.X_SR_LATCH.nand_0.drain_mna VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X37 VGND.t49 X_TIMER.qb_sr X_TIMER.q_sr VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X38 uo_out[0].t3 X_TIMER.out_inv1 VGND.t46 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X39 X_TIMER.out_inv3 uo_out[0].t10 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X40 X_TIMER.X_COMP_P_BOTTOM.tail.t1 X_TIMER.v0p6 X_TIMER.X_COMP_P_BOTTOM.latch_right.t1 VPWR.t1 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X41 uo_out[0].t0 X_TIMER.out_inv1 VGND.t45 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X42 VGND.t50 X_TIMER.X_COMP_P_TOP.latch_right.t7 X_TIMER.X_SR_LATCH.IN_R.t1 VGND.t34 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
X43 VGND.t12 X_TIMER.X_COMP_P_TOP.latch_left.t4 X_TIMER.X_COMP_P_TOP.latch_left.t5 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X44 ua[2].t4 X_TIMER.out_inv3 VGND.t25 VGND.t24 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.35
X45 X_TIMER.qb_sr X_TIMER.X_SR_LATCH.IN_S.t3 a_1347_2994# VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X46 X_TIMER.X_COMP_P_BOTTOM.tail.t0 X_TIMER.v0p6 X_TIMER.X_COMP_P_BOTTOM.latch_right.t0 VPWR.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X47 VGND.t14 X_TIMER.q_sr X_TIMER.qb_sr VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X48 X_TIMER.X_COMP_P_TOP.latch_right.t4 ua[0].t2 X_TIMER.X_COMP_P_TOP.tail.t5 VPWR.t11 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X49 VGND.t23 X_TIMER.out_inv3 ua[2].t3 VGND.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X50 VPWR.t20 X_TIMER.X_COMP_P_BOTTOM.out_left.t0 X_TIMER.X_COMP_P_BOTTOM.out_left.t1 VPWR.t19 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
X51 VPWR.t42 X_TIMER.X_SR_LATCH.nand_0.IN_A X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B VPWR.t41 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X52 VGND.t21 X_TIMER.out_inv3 ua[2].t2 VGND.t20 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X53 X_TIMER.X_COMP_P_BOTTOM.tail.t4 ua[1].t2 X_TIMER.X_COMP_P_BOTTOM.latch_left.t4 VPWR.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X54 X_TIMER.bias_3 X_TIMER.bias_2 VGND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=7
X55 X_TIMER.bias_1 X_TIMER.bias_p VGND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=7
X56 ua[2].t1 X_TIMER.out_inv3 VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8_lvt ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.35
X57 ua[2].t0 X_TIMER.out_inv3 VGND.t17 VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X58 X_TIMER.X_COMP_P_BOTTOM.tail.t5 ua[1].t3 X_TIMER.X_COMP_P_BOTTOM.latch_left.t3 VPWR.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X59 X_TIMER.X_COMP_P_TOP.out_left.t1 X_TIMER.X_COMP_P_TOP.out_left.t0 VPWR.t40 VPWR.t39 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
X60 X_TIMER.X_COMP_P_BOTTOM.latch_left.t2 X_TIMER.X_COMP_P_BOTTOM.latch_left.t1 VGND.t38 VGND.t37 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X61 X_TIMER.X_SR_LATCH.nand_0.IN_A X_TIMER.X_SR_LATCH.IN_R.t3 VGND.t47 VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X62 X_TIMER.v1p2 VPWR VGND.t39 sky130_fd_pr__res_xhigh_po_1p41 l=7
X63 X_TIMER.bias_3 X_TIMER.bias_n VGND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=7
X64 VGND.t10 X_TIMER.X_COMP_P_TOP.latch_left.t8 X_TIMER.X_COMP_P_TOP.latch_right.t0 VGND.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
X65 VGND.t27 X_TIMER.X_COMP_P_TOP.latch_right.t1 X_TIMER.X_COMP_P_TOP.latch_right.t2 VGND.t26 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X66 a_1723_2994# X_TIMER.qb_sr VPWR.t44 VPWR.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X67 X_TIMER.X_SR_LATCH.nand_0.drain_mna X_TIMER.X_SR_LATCH.nand_0.IN_A VGND.t48 VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X68 X_TIMER.X_COMP_P_BOTTOM.out_left.t2 X_TIMER.X_COMP_P_BOTTOM.latch_left.t7 VGND.t36 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
X69 X_TIMER.X_COMP_P_TOP.latch_left.t0 X_TIMER.v1p2 X_TIMER.X_COMP_P_TOP.tail.t2 VPWR.t12 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X70 a_1347_2994# X_TIMER.q_sr VPWR.t16 VPWR.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X71 X_TIMER.q_sr X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B VGND.t8 VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X72 VGND.t35 X_TIMER.X_COMP_P_TOP.latch_right.t8 X_TIMER.X_COMP_P_TOP.latch_left.t6 VGND.t34 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
X73 X_TIMER.X_COMP_P_TOP.latch_right.t3 ua[0].t3 X_TIMER.X_COMP_P_TOP.tail.t7 VPWR.t12 sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X74 X_TIMER.out_inv3 uo_out[0].t11 VPWR.t3 VPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X75 X_TIMER.X_COMP_P_BOTTOM.latch_right.t4 X_TIMER.X_COMP_P_BOTTOM.latch_left.t8 VGND.t6 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
R0 uo_out[0].n6 uo_out[0].t5 411.07
R1 uo_out[0].n5 uo_out[0].t9 411.07
R2 uo_out[0].n4 uo_out[0].t10 411.07
R3 uo_out[0].n3 uo_out[0].t6 411.07
R4 uo_out[0].n6 uo_out[0].t11 400.375
R5 uo_out[0].n5 uo_out[0].t7 400.375
R6 uo_out[0].n4 uo_out[0].t8 400.375
R7 uo_out[0].n2 uo_out[0].t4 395.873
R8 uo_out[0].n1 uo_out[0].t1 228.959
R9 uo_out[0].n0 uo_out[0].t2 228.959
R10 uo_out[0].n1 uo_out[0].t3 84.8864
R11 uo_out[0].n0 uo_out[0].t0 84.8864
R12 uo_out[0].n7 uo_out[0] 39.2126
R13 uo_out[0] uo_out[0].n6 28.1147
R14 uo_out[0].n3 uo_out[0].n2 4.50234
R15 uo_out[0].n1 uo_out[0] 0.8755
R16 uo_out[0].n2 uo_out[0] 0.800132
R17 uo_out[0] uo_out[0].n3 0.382853
R18 uo_out[0] uo_out[0].n4 0.382853
R19 uo_out[0] uo_out[0].n5 0.382853
R20 uo_out[0].n3 uo_out[0] 0.378389
R21 uo_out[0].n4 uo_out[0] 0.378389
R22 uo_out[0].n5 uo_out[0] 0.378389
R23 uo_out[0].n6 uo_out[0] 0.378389
R24 uo_out[0].n7 uo_out[0] 0.120692
R25 uo_out[0] uo_out[0].n7 0.116241
R26 uo_out[0] uo_out[0].n1 0.0924118
R27 uo_out[0] uo_out[0].n0 0.0924118
R28 VPWR.n92 VPWR.n41 5809.41
R29 VPWR.n92 VPWR.n91 5809.41
R30 VPWR.n100 VPWR.n36 5809.41
R31 VPWR.n100 VPWR.n99 5809.41
R32 VPWR.n87 VPWR.n43 5784.71
R33 VPWR.n89 VPWR.n43 5784.71
R34 VPWR.n69 VPWR.n67 5784.71
R35 VPWR.n69 VPWR.n68 5784.71
R36 VPWR.n121 VPWR.n117 4912.94
R37 VPWR.n118 VPWR.n115 4912.94
R38 VPWR.n59 VPWR.n38 4912.94
R39 VPWR.n96 VPWR.n38 4912.94
R40 VPWR.n59 VPWR.n23 4912.94
R41 VPWR.n96 VPWR.n23 4912.94
R42 VPWR.n153 VPWR.n6 4912.94
R43 VPWR.n152 VPWR.n6 4912.94
R44 VPWR.n152 VPWR.n5 4912.94
R45 VPWR.n153 VPWR.n5 4912.94
R46 VPWR.n104 VPWR.n32 4208.75
R47 VPWR.n108 VPWR.n107 4207.06
R48 VPWR.n75 VPWR.n65 4207.06
R49 VPWR.n78 VPWR.n57 4205.22
R50 VPWR.n87 VPWR.n47 4020
R51 VPWR.n90 VPWR.n89 4020
R52 VPWR.n67 VPWR.n11 4020
R53 VPWR.n68 VPWR.n12 4020
R54 VPWR.n47 VPWR.n41 3998.82
R55 VPWR.n91 VPWR.n90 3998.82
R56 VPWR.n36 VPWR.n11 3998.82
R57 VPWR.n99 VPWR.n12 3998.82
R58 VPWR.n57 VPWR.n26 3409.41
R59 VPWR.n108 VPWR.n26 3409.41
R60 VPWR.n65 VPWR.n14 3409.41
R61 VPWR.n32 VPWR.n14 3409.41
R62 VPWR.n47 VPWR.n42 1789.41
R63 VPWR.n90 VPWR.n42 1789.41
R64 VPWR.n148 VPWR.n11 1789.41
R65 VPWR.n148 VPWR.n12 1789.41
R66 VPWR.n119 VPWR.n118 1373.18
R67 VPWR.n121 VPWR.n120 1373.18
R68 VPWR.n194 VPWR.n181 1297.82
R69 VPWR.n194 VPWR.n162 1289.14
R70 VPWR.n197 VPWR.n162 1146.76
R71 VPWR.n187 VPWR.n181 1136.47
R72 VPWR.n61 VPWR.n56 981.356
R73 VPWR.n64 VPWR.n63 981.356
R74 VPWR.n51 VPWR.n13 981.356
R75 VPWR.n50 VPWR.n27 981.356
R76 VPWR.n168 VPWR.n167 928.236
R77 VPWR.n168 VPWR.n163 928.236
R78 VPWR.n179 VPWR.n163 928.236
R79 VPWR.n180 VPWR.n179 928.236
R80 VPWR.n180 VPWR.n160 928.236
R81 VPWR.n197 VPWR.n160 924.707
R82 VPWR.n78 VPWR.n56 801.5
R83 VPWR.n104 VPWR.n27 800.322
R84 VPWR.n62 VPWR.n26 797.648
R85 VPWR.n63 VPWR.n62 797.648
R86 VPWR.n75 VPWR.n56 797.648
R87 VPWR.n146 VPWR.n13 797.648
R88 VPWR.n146 VPWR.n14 797.648
R89 VPWR.n107 VPWR.n27 797.648
R90 VPWR.n116 VPWR.n114 524.048
R91 VPWR.n123 VPWR.n114 524.048
R92 VPWR.n122 VPWR.n116 524.048
R93 VPWR.n123 VPWR.n122 524.048
R94 VPWR.n93 VPWR.n40 447.06
R95 VPWR.n101 VPWR.n34 447.06
R96 VPWR.n70 VPWR.n66 444.515
R97 VPWR.n86 VPWR.n81 444.515
R98 VPWR.n66 VPWR.n10 428.8
R99 VPWR.n86 VPWR.n85 428.8
R100 VPWR.n34 VPWR.n10 426.541
R101 VPWR.n85 VPWR.n40 426.541
R102 VPWR.t17 VPWR.t10 417.711
R103 VPWR.t43 VPWR.t27 417.711
R104 VPWR.t23 VPWR.t15 411.909
R105 VPWR.t13 VPWR.t41 397.406
R106 VPWR.t6 VPWR.t2 381.45
R107 VPWR.t6 VPWR.t4 381.45
R108 VPWR.t4 VPWR.t8 381.45
R109 VPWR.t31 VPWR.t8 381.45
R110 VPWR.t29 VPWR.t31 381.45
R111 VPWR.t17 VPWR.t29 380
R112 VPWR.n144 VPWR.n15 363.671
R113 VPWR.n55 VPWR.n54 363.671
R114 VPWR.n143 VPWR.n16 363.295
R115 VPWR.n53 VPWR.n52 363.295
R116 VPWR.n74 VPWR.n15 362.37
R117 VPWR.n79 VPWR.n55 362.37
R118 VPWR.n103 VPWR.n16 361.584
R119 VPWR.n52 VPWR.n28 361.584
R120 VPWR.n158 VPWR.t30 228.663
R121 VPWR.n182 VPWR.t18 228.663
R122 VPWR.n185 VPWR.t14 228.663
R123 VPWR.n165 VPWR.t3 228.663
R124 VPWR.n171 VPWR.t7 228.663
R125 VPWR.n173 VPWR.t5 228.663
R126 VPWR.n176 VPWR.t9 228.663
R127 VPWR.n174 VPWR.t32 228.663
R128 VPWR.n190 VPWR.n189 202.965
R129 VPWR.n150 VPWR.n149 190.871
R130 VPWR.n149 VPWR.n10 190.871
R131 VPWR.n85 VPWR.n84 190.871
R132 VPWR.n84 VPWR.n83 190.871
R133 VPWR.n147 VPWR.t39 175.422
R134 VPWR.t25 VPWR.t37 171.423
R135 VPWR.n106 VPWR.n29 143.065
R136 VPWR.n76 VPWR.n60 135.065
R137 VPWR.n192 VPWR.t16 114.451
R138 VPWR.n184 VPWR.t44 114.451
R139 VPWR.n169 VPWR.n166 99.0123
R140 VPWR.n169 VPWR.n164 99.0123
R141 VPWR.n178 VPWR.n164 99.0123
R142 VPWR.n178 VPWR.n159 99.0123
R143 VPWR.n199 VPWR.n159 99.0123
R144 VPWR.n199 VPWR.n198 98.6358
R145 VPWR.n188 VPWR.n187 97.1505
R146 VPWR.n187 VPWR.t13 92.5005
R147 VPWR.n167 VPWR.n166 92.5005
R148 VPWR.t2 VPWR.n167 92.5005
R149 VPWR.n169 VPWR.n168 92.5005
R150 VPWR.n168 VPWR.t6 92.5005
R151 VPWR.n164 VPWR.n163 92.5005
R152 VPWR.t4 VPWR.n163 92.5005
R153 VPWR.n179 VPWR.n178 92.5005
R154 VPWR.n179 VPWR.t8 92.5005
R155 VPWR.n180 VPWR.n159 92.5005
R156 VPWR.t31 VPWR.n180 92.5005
R157 VPWR.n199 VPWR.n160 92.5005
R158 VPWR.t29 VPWR.n160 92.5005
R159 VPWR.n198 VPWR.n197 92.5005
R160 VPWR.n197 VPWR.t17 92.5005
R161 VPWR.n145 VPWR.n144 85.0829
R162 VPWR.n145 VPWR.n4 85.0829
R163 VPWR.n110 VPWR.n24 85.0829
R164 VPWR.n54 VPWR.n24 85.0829
R165 VPWR.t41 VPWR.n186 69.6188
R166 VPWR.n196 VPWR.t43 68.1684
R167 VPWR.n195 VPWR.t15 68.1684
R168 VPWR.n150 VPWR.n9 66.7857
R169 VPWR.n83 VPWR.n25 66.7857
R170 VPWR.n151 VPWR.n8 66.1931
R171 VPWR.n82 VPWR.n44 66.1931
R172 VPWR.n105 VPWR.n30 61.6251
R173 VPWR.n77 VPWR.n58 61.4433
R174 VPWR.t10 VPWR.n196 59.4661
R175 VPWR.t27 VPWR.n195 59.4661
R176 VPWR.n186 VPWR.t23 58.0158
R177 VPWR.n31 VPWR.n4 52.3937
R178 VPWR.n110 VPWR.n109 52.3937
R179 VPWR.n154 VPWR.n3 51.2005
R180 VPWR.n111 VPWR.n22 51.2005
R181 VPWR.n183 VPWR.n162 49.3505
R182 VPWR.n194 VPWR.n193 49.3505
R183 VPWR.n190 VPWR.n181 46.2505
R184 VPWR.n186 VPWR.n181 46.2505
R185 VPWR.n196 VPWR.n162 46.2505
R186 VPWR.n195 VPWR.n194 46.2505
R187 VPWR.n118 VPWR.n114 37.0005
R188 VPWR.n122 VPWR.n121 37.0005
R189 VPWR.n75 VPWR.n74 37.0005
R190 VPWR.n76 VPWR.n75 37.0005
R191 VPWR.n72 VPWR.n5 37.0005
R192 VPWR.n45 VPWR.n5 37.0005
R193 VPWR.n33 VPWR.n6 37.0005
R194 VPWR.n29 VPWR.n6 37.0005
R195 VPWR.n104 VPWR.n103 37.0005
R196 VPWR.n105 VPWR.n104 37.0005
R197 VPWR.n146 VPWR.n145 37.0005
R198 VPWR.n147 VPWR.n146 37.0005
R199 VPWR.n107 VPWR.n28 37.0005
R200 VPWR.n107 VPWR.n106 37.0005
R201 VPWR.n96 VPWR.n95 37.0005
R202 VPWR.n97 VPWR.n96 37.0005
R203 VPWR.n59 VPWR.n49 37.0005
R204 VPWR.n60 VPWR.n59 37.0005
R205 VPWR.n79 VPWR.n78 37.0005
R206 VPWR.n78 VPWR.n77 37.0005
R207 VPWR.n62 VPWR.n24 37.0005
R208 VPWR.n62 VPWR.n7 37.0005
R209 VPWR.t21 VPWR.t1 30.5401
R210 VPWR.t19 VPWR.n37 30.1765
R211 VPWR.n130 VPWR.t22 29.4286
R212 VPWR.n129 VPWR.t26 29.4286
R213 VPWR.n139 VPWR.t40 29.4286
R214 VPWR.n138 VPWR.t20 29.4286
R215 VPWR.n73 VPWR.n70 26.6787
R216 VPWR.n81 VPWR.n80 26.6787
R217 VPWR.n94 VPWR.n93 26.63
R218 VPWR.n102 VPWR.n101 26.63
R219 VPWR.n124 VPWR.t34 23.3739
R220 VPWR.n111 VPWR.t38 23.0294
R221 VPWR.n154 VPWR.t36 23.0294
R222 VPWR.n48 VPWR.n22 19.0689
R223 VPWR.n71 VPWR.n3 19.0689
R224 VPWR.n102 VPWR.n33 17.4344
R225 VPWR.n95 VPWR.n94 17.4344
R226 VPWR.n109 VPWR.n25 16.8923
R227 VPWR.n31 VPWR.n9 16.8923
R228 VPWR.n73 VPWR.n72 16.6793
R229 VPWR.n80 VPWR.n49 16.6793
R230 VPWR.n58 VPWR.n43 14.4131
R231 VPWR.n100 VPWR.n30 14.4131
R232 VPWR.n189 VPWR.t24 14.283
R233 VPWR.n189 VPWR.t42 14.283
R234 VPWR.n93 VPWR.n92 14.2313
R235 VPWR.n92 VPWR.n30 14.2313
R236 VPWR.n70 VPWR.n69 14.2313
R237 VPWR.n69 VPWR.n58 14.2313
R238 VPWR.n149 VPWR.n148 14.2313
R239 VPWR.n148 VPWR.n147 14.2313
R240 VPWR.n101 VPWR.n100 14.2313
R241 VPWR.n84 VPWR.n42 14.2313
R242 VPWR.n42 VPWR.n7 14.2313
R243 VPWR.n81 VPWR.n43 14.2313
R244 VPWR.n88 VPWR.n45 8.7261
R245 VPWR.n32 VPWR.n31 7.11588
R246 VPWR.t19 VPWR.n32 7.11588
R247 VPWR.n65 VPWR.n3 7.11588
R248 VPWR.n65 VPWR.t25 7.11588
R249 VPWR.n50 VPWR.n16 7.11588
R250 VPWR.n50 VPWR.t19 7.11588
R251 VPWR.n64 VPWR.n15 7.11588
R252 VPWR.t25 VPWR.n64 7.11588
R253 VPWR.n61 VPWR.n55 7.11588
R254 VPWR.n61 VPWR.t21 7.11588
R255 VPWR.n52 VPWR.n51 7.11588
R256 VPWR.n51 VPWR.t39 7.11588
R257 VPWR.n57 VPWR.n22 7.11588
R258 VPWR.t21 VPWR.n57 7.11588
R259 VPWR.n109 VPWR.n108 7.11588
R260 VPWR.n108 VPWR.t39 7.11588
R261 VPWR.n117 VPWR.n116 5.78175
R262 VPWR.n123 VPWR.n115 5.78175
R263 VPWR.n154 VPWR.n153 5.78175
R264 VPWR.n153 VPWR.t35 5.78175
R265 VPWR.n67 VPWR.n8 5.78175
R266 VPWR.n67 VPWR.n46 5.78175
R267 VPWR.n152 VPWR.n151 5.78175
R268 VPWR.t35 VPWR.n152 5.78175
R269 VPWR.n99 VPWR.n34 5.78175
R270 VPWR.n99 VPWR.n98 5.78175
R271 VPWR.n68 VPWR.n66 5.78175
R272 VPWR.n68 VPWR.n46 5.78175
R273 VPWR.n36 VPWR.n35 5.78175
R274 VPWR.n98 VPWR.n36 5.78175
R275 VPWR.n91 VPWR.n39 5.78175
R276 VPWR.n91 VPWR.n37 5.78175
R277 VPWR.n82 VPWR.n38 5.78175
R278 VPWR.n38 VPWR.t37 5.78175
R279 VPWR.n89 VPWR.n44 5.78175
R280 VPWR.n89 VPWR.n88 5.78175
R281 VPWR.n87 VPWR.n86 5.78175
R282 VPWR.n88 VPWR.n87 5.78175
R283 VPWR.n41 VPWR.n40 5.78175
R284 VPWR.n41 VPWR.n37 5.78175
R285 VPWR.n111 VPWR.n23 5.78175
R286 VPWR.n23 VPWR.t37 5.78175
R287 VPWR.n166 VPWR.n165 4.74533
R288 VPWR.n103 VPWR.n102 4.7119
R289 VPWR.n94 VPWR.n28 4.7119
R290 VPWR.n74 VPWR.n73 4.70083
R291 VPWR.n80 VPWR.n79 4.70083
R292 VPWR.n200 VPWR.n199 4.6505
R293 VPWR.n198 VPWR.n161 4.6505
R294 VPWR.n170 VPWR.n169 4.6505
R295 VPWR.n172 VPWR.n164 4.6505
R296 VPWR.n178 VPWR.n177 4.6505
R297 VPWR.n175 VPWR.n159 4.6505
R298 VPWR.n119 VPWR.n117 4.16148
R299 VPWR.n120 VPWR.n115 4.16148
R300 VPWR.n132 VPWR 4.11685
R301 VPWR.t35 VPWR.n7 3.81795
R302 VPWR.n134 VPWR.n133 3.36117
R303 VPWR.n191 VPWR.n190 3.1005
R304 VPWR.n113 VPWR.n112 2.9268
R305 VPWR.n155 VPWR.n1 2.92408
R306 VPWR.n156 VPWR.n155 2.92408
R307 VPWR.n112 VPWR.n21 2.92137
R308 VPWR.n141 VPWR 2.25915
R309 VPWR.n131 VPWR 2.19312
R310 VPWR.n71 VPWR.n8 1.77828
R311 VPWR.n48 VPWR.n44 1.77828
R312 VPWR.n120 VPWR.t33 1.61687
R313 VPWR.t33 VPWR.n119 1.61687
R314 VPWR.n151 VPWR.n150 1.3042
R315 VPWR.n83 VPWR.n82 1.3042
R316 VPWR.n140 VPWR 1.20337
R317 VPWR.n154 VPWR.n4 1.19372
R318 VPWR.n111 VPWR.n110 1.19372
R319 VPWR.t0 VPWR.n97 1.0912
R320 VPWR.n64 VPWR.n61 1.01745
R321 VPWR.n63 VPWR.n13 1.01745
R322 VPWR.n51 VPWR.n50 1.01745
R323 VPWR.n19 VPWR 0.941142
R324 VPWR.n133 VPWR 0.856789
R325 VPWR.n20 VPWR.n0 0.830381
R326 VPWR VPWR.n191 0.66955
R327 VPWR.n203 VPWR 0.662254
R328 VPWR.n135 VPWR 0.590885
R329 VPWR.n183 VPWR 0.568535
R330 VPWR.n193 VPWR 0.564096
R331 VPWR VPWR.n188 0.55213
R332 VPWR.t12 VPWR.n46 0.54585
R333 VPWR.n98 VPWR.t11 0.54585
R334 VPWR.n203 VPWR.n202 0.424031
R335 VPWR.n170 VPWR 0.417194
R336 VPWR.n172 VPWR 0.417194
R337 VPWR.n177 VPWR 0.417194
R338 VPWR VPWR.n175 0.417194
R339 VPWR.n202 VPWR.n157 0.416109
R340 VPWR.n161 VPWR 0.41479
R341 VPWR.n136 VPWR 0.395992
R342 VPWR.n144 VPWR.n143 0.376971
R343 VPWR.n54 VPWR.n53 0.376971
R344 VPWR.n126 VPWR.n125 0.371147
R345 VPWR.n201 VPWR.n200 0.352871
R346 VPWR.n155 VPWR.n154 0.344944
R347 VPWR.n112 VPWR.n111 0.344944
R348 VPWR.n191 VPWR 0.32387
R349 VPWR.n124 VPWR.n123 0.3105
R350 VPWR.n72 VPWR.n71 0.307571
R351 VPWR.n49 VPWR.n48 0.307571
R352 VPWR.n140 VPWR.n139 0.27529
R353 VPWR.n138 VPWR.n137 0.27529
R354 VPWR.n131 VPWR.n130 0.27529
R355 VPWR.n137 VPWR 0.270402
R356 VPWR.n125 VPWR.n124 0.259149
R357 VPWR.n128 VPWR.n127 0.234786
R358 VPWR.n202 VPWR.n201 0.225984
R359 VPWR.n21 VPWR.n20 0.209875
R360 VPWR.n157 VPWR.n156 0.209435
R361 VPWR.n184 VPWR.n183 0.202254
R362 VPWR.n193 VPWR.n192 0.202254
R363 VPWR.n77 VPWR.n76 0.182283
R364 VPWR.n60 VPWR.n45 0.182283
R365 VPWR.n88 VPWR.n46 0.182283
R366 VPWR.t1 VPWR.t12 0.182283
R367 VPWR.t25 VPWR.t21 0.182283
R368 VPWR.t35 VPWR.t37 0.182283
R369 VPWR.n147 VPWR.n7 0.182283
R370 VPWR.t19 VPWR.t39 0.182283
R371 VPWR.n98 VPWR.n37 0.182283
R372 VPWR.t11 VPWR.t0 0.182283
R373 VPWR.n97 VPWR.n29 0.182283
R374 VPWR.n106 VPWR.n105 0.182283
R375 VPWR.n35 VPWR.n33 0.178728
R376 VPWR.n95 VPWR.n39 0.178728
R377 VPWR.n129 VPWR.n128 0.177874
R378 VPWR.n142 VPWR.n141 0.169731
R379 VPWR.n19 VPWR.n17 0.162038
R380 VPWR.n136 VPWR.n135 0.152423
R381 VPWR.n133 VPWR.n132 0.152423
R382 VPWR.n143 VPWR.n142 0.133357
R383 VPWR.n53 VPWR.n17 0.133357
R384 VPWR.n125 VPWR.n0 0.122632
R385 VPWR.n188 VPWR.n185 0.120065
R386 VPWR.n127 VPWR.n126 0.116433
R387 VPWR.n128 VPWR.n19 0.101757
R388 VPWR.n35 VPWR.n9 0.0977152
R389 VPWR.n39 VPWR.n25 0.0977152
R390 VPWR.n185 VPWR 0.0956087
R391 VPWR.n200 VPWR.n158 0.0953276
R392 VPWR.n182 VPWR.n161 0.0953276
R393 VPWR.n171 VPWR.n170 0.0953276
R394 VPWR.n173 VPWR.n172 0.0953276
R395 VPWR.n177 VPWR.n176 0.0953276
R396 VPWR.n175 VPWR.n174 0.0953276
R397 VPWR.n134 VPWR.n18 0.0882225
R398 VPWR VPWR.n158 0.075931
R399 VPWR VPWR.n182 0.075931
R400 VPWR.n165 VPWR 0.075931
R401 VPWR VPWR.n171 0.075931
R402 VPWR VPWR.n173 0.075931
R403 VPWR.n176 VPWR 0.075931
R404 VPWR.n174 VPWR 0.075931
R405 VPWR.n113 VPWR.n20 0.068875
R406 VPWR.n157 VPWR.n1 0.067875
R407 VPWR.n156 VPWR.n2 0.0652508
R408 VPWR.n201 VPWR 0.0648236
R409 VPWR.n126 VPWR.n1 0.06425
R410 VPWR.n21 VPWR.n2 0.0640173
R411 VPWR.n126 VPWR.n113 0.064
R412 VPWR VPWR.n203 0.061493
R413 VPWR VPWR.n184 0.0597105
R414 VPWR.n192 VPWR 0.0597105
R415 VPWR.n135 VPWR.n134 0.0323455
R416 VPWR.n127 VPWR.n2 0.0187405
R417 VPWR.n203 VPWR.n0 0.0120348
R418 VPWR.n142 VPWR.n17 0.00146154
R419 VPWR.n18 VPWR 0.00119261
R420 VPWR.n141 VPWR.n140 0.0010123
R421 VPWR.n137 VPWR.n136 0.0010123
R422 VPWR.n132 VPWR.n131 0.0010123
R423 VPWR.n18 VPWR 0.00100029
R424 VPWR.n139 VPWR.n138 0.000849162
R425 VPWR.n130 VPWR.n129 0.000849162
R426 X_TIMER.X_COMP_P_BOTTOM.latch_right.n4 X_TIMER.X_COMP_P_BOTTOM.latch_right.t7 114.778
R427 X_TIMER.X_COMP_P_BOTTOM.latch_right.n4 X_TIMER.X_COMP_P_BOTTOM.latch_right.t8 106.572
R428 X_TIMER.X_COMP_P_BOTTOM.latch_right.n3 X_TIMER.X_COMP_P_BOTTOM.latch_right.t1 28.4736
R429 X_TIMER.X_COMP_P_BOTTOM.latch_right.n3 X_TIMER.X_COMP_P_BOTTOM.latch_right.t3 28.057
R430 X_TIMER.X_COMP_P_BOTTOM.latch_right.n0 X_TIMER.X_COMP_P_BOTTOM.latch_right.t0 27.8467
R431 X_TIMER.X_COMP_P_BOTTOM.latch_right.n0 X_TIMER.X_COMP_P_BOTTOM.latch_right.t2 27.4301
R432 X_TIMER.X_COMP_P_BOTTOM.latch_right.n1 X_TIMER.X_COMP_P_BOTTOM.latch_right.t6 22.0141
R433 X_TIMER.X_COMP_P_BOTTOM.latch_right.n0 X_TIMER.X_COMP_P_BOTTOM.latch_right.t4 20.4334
R434 X_TIMER.X_COMP_P_BOTTOM.latch_right.n2 X_TIMER.X_COMP_P_BOTTOM.latch_right.n1 0.582966
R435 X_TIMER.X_COMP_P_BOTTOM.latch_right.n2 X_TIMER.X_COMP_P_BOTTOM.latch_right.n4 1.69623
R436 X_TIMER.X_COMP_P_BOTTOM.latch_right.n2 X_TIMER.X_COMP_P_BOTTOM.latch_right.t5 95.1763
R437 X_TIMER.X_COMP_P_BOTTOM.latch_right X_TIMER.X_COMP_P_BOTTOM.latch_right.n0 14.0375
R438 X_TIMER.X_COMP_P_BOTTOM.latch_right X_TIMER.X_COMP_P_BOTTOM.latch_right.n1 0.612947
R439 X_TIMER.X_COMP_P_BOTTOM.latch_right X_TIMER.X_COMP_P_BOTTOM.latch_right.n3 0.516125
R440 VGND.n133 VGND.n132 5.73231e+06
R441 VGND.n256 VGND.n255 3.08487e+06
R442 VGND.n255 VGND.n254 11223.8
R443 VGND.n215 VGND.n68 9119.94
R444 VGND.n216 VGND.n68 9119.94
R445 VGND.n215 VGND.n69 9119.94
R446 VGND.n216 VGND.n69 9119.94
R447 VGND.n248 VGND.n227 8494.18
R448 VGND.n248 VGND.n238 8494.18
R449 VGND.n253 VGND.n228 8494.18
R450 VGND.n234 VGND.n228 8494.18
R451 VGND.n37 VGND.n27 8494.18
R452 VGND.n257 VGND.n27 8494.18
R453 VGND.n275 VGND.n21 8494.18
R454 VGND.n275 VGND.n26 8494.18
R455 VGND.n274 VGND.n34 7555.55
R456 VGND.n237 VGND.n236 7120.97
R457 VGND.n240 VGND.n237 7120.97
R458 VGND.n249 VGND.n229 7120.97
R459 VGND.n249 VGND.n235 7120.97
R460 VGND.n36 VGND.n31 7120.97
R461 VGND.n47 VGND.n31 7120.97
R462 VGND.n39 VGND.n32 7120.97
R463 VGND.n46 VGND.n32 7120.97
R464 VGND.n38 VGND.n33 7120.97
R465 VGND.n258 VGND.n33 7120.97
R466 VGND.n160 VGND.n80 5440.68
R467 VGND.n299 VGND.n7 5440.68
R468 VGND.n280 VGND.n22 5440.68
R469 VGND.n280 VGND.n23 5440.68
R470 VGND.n138 VGND.n96 5255.26
R471 VGND.n124 VGND.n120 5255.26
R472 VGND.n29 VGND.n22 5255.26
R473 VGND.n29 VGND.n23 5255.26
R474 VGND.n134 VGND.n100 4536.79
R475 VGND.n135 VGND.n100 4536.79
R476 VGND.n181 VGND.n71 4536.79
R477 VGND.n181 VGND.n72 4536.79
R478 VGND.n291 VGND.n19 4536.79
R479 VGND.n292 VGND.n19 4536.79
R480 VGND.n131 VGND.n102 4536.79
R481 VGND.n131 VGND.n101 4536.79
R482 VGND.n96 VGND.n79 4131.21
R483 VGND.n146 VGND.n84 4131.21
R484 VGND.n159 VGND.n85 4131.21
R485 VGND.n148 VGND.n147 4131.21
R486 VGND.n154 VGND.n83 4131.21
R487 VGND.n120 VGND.n6 4131.21
R488 VGND.n113 VGND.n112 4131.21
R489 VGND.n293 VGND.n10 4131.21
R490 VGND.n119 VGND.n11 4131.21
R491 VGND.n298 VGND.n12 4131.21
R492 VGND.n160 VGND.n79 3945.79
R493 VGND.n146 VGND.n97 3945.79
R494 VGND.n159 VGND.n84 3945.79
R495 VGND.n147 VGND.n94 3945.79
R496 VGND.n148 VGND.n83 3945.79
R497 VGND.n299 VGND.n6 3945.79
R498 VGND.n113 VGND.n107 3945.79
R499 VGND.n112 VGND.n10 3945.79
R500 VGND.n119 VGND.n106 3945.79
R501 VGND.n298 VGND.n11 3945.79
R502 VGND.n264 VGND.n256 3787.12
R503 VGND.n134 VGND.n97 3227.32
R504 VGND.n85 VGND.n71 3227.32
R505 VGND.n135 VGND.n94 3227.32
R506 VGND.n154 VGND.n72 3227.32
R507 VGND.n107 VGND.n102 3227.32
R508 VGND.n293 VGND.n292 3227.32
R509 VGND.n106 VGND.n101 3227.32
R510 VGND.n291 VGND.n12 3227.32
R511 VGND.t33 VGND.n274 3048.25
R512 VGND.n264 VGND.n48 2152.87
R513 VGND.n61 VGND.n52 2131.24
R514 VGND.n254 VGND.n226 2128.64
R515 VGND.n221 VGND.n53 1904.94
R516 VGND.n225 VGND.n49 1692.69
R517 VGND.n211 VGND.n209 1523.85
R518 VGND.n209 VGND.n208 1523.85
R519 VGND.n205 VGND.n204 1523.85
R520 VGND.n236 VGND.n227 1373.21
R521 VGND.n241 VGND.n235 1373.21
R522 VGND.n241 VGND.n240 1373.21
R523 VGND.n240 VGND.n238 1373.21
R524 VGND.n253 VGND.n229 1373.21
R525 VGND.n229 VGND.n224 1373.21
R526 VGND.n236 VGND.n224 1373.21
R527 VGND.n235 VGND.n234 1373.21
R528 VGND.n37 VGND.n36 1373.21
R529 VGND.n265 VGND.n46 1373.21
R530 VGND.n265 VGND.n47 1373.21
R531 VGND.n257 VGND.n47 1373.21
R532 VGND.n273 VGND.n38 1373.21
R533 VGND.n273 VGND.n39 1373.21
R534 VGND.n39 VGND.n35 1373.21
R535 VGND.n36 VGND.n35 1373.21
R536 VGND.n258 VGND.n26 1373.21
R537 VGND.n263 VGND.n258 1373.21
R538 VGND.n263 VGND.n46 1373.21
R539 VGND.n38 VGND.n21 1373.21
R540 VGND.n256 VGND.n49 1351.14
R541 VGND.n138 VGND.n94 1309.47
R542 VGND.n148 VGND.n93 1309.47
R543 VGND.n93 VGND.n79 1309.47
R544 VGND.n154 VGND.n80 1309.47
R545 VGND.n155 VGND.n85 1309.47
R546 VGND.n155 VGND.n154 1309.47
R547 VGND.n149 VGND.n84 1309.47
R548 VGND.n149 VGND.n148 1309.47
R549 VGND.n142 VGND.n97 1309.47
R550 VGND.n142 VGND.n94 1309.47
R551 VGND.n13 VGND.n6 1309.47
R552 VGND.n13 VGND.n11 1309.47
R553 VGND.n124 VGND.n106 1309.47
R554 VGND.n12 VGND.n7 1309.47
R555 VGND.n126 VGND.n106 1309.47
R556 VGND.n126 VGND.n107 1309.47
R557 VGND.n111 VGND.n11 1309.47
R558 VGND.n112 VGND.n111 1309.47
R559 VGND.n294 VGND.n12 1309.47
R560 VGND.n294 VGND.n293 1309.47
R561 VGND.t28 VGND.n81 1288.91
R562 VGND.t5 VGND.n82 1288.91
R563 VGND.t28 VGND.n95 1231.06
R564 VGND.t5 VGND.n81 1231.06
R565 VGND.t31 VGND.n133 1006.9
R566 VGND.t31 VGND.n95 1006.9
R567 VGND.n82 VGND.t37 1006.9
R568 VGND.n182 VGND.t37 1006.9
R569 VGND.n214 VGND.n67 592.566
R570 VGND.n247 VGND.n239 551.907
R571 VGND.n247 VGND.n246 551.907
R572 VGND.n252 VGND.n230 551.907
R573 VGND.n233 VGND.n230 551.907
R574 VGND.n44 VGND.n43 551.907
R575 VGND.n43 VGND.n42 551.907
R576 VGND.n217 VGND.n67 546.303
R577 VGND.n169 VGND.n50 528.745
R578 VGND.n260 VGND.n25 528.566
R579 VGND.n210 VGND.n184 503.861
R580 VGND.n244 VGND.n243 462.683
R581 VGND.n245 VGND.n244 462.683
R582 VGND.n251 VGND.n250 462.683
R583 VGND.n250 VGND.n232 462.683
R584 VGND.n271 VGND.n41 462.683
R585 VGND.n45 VGND.n41 462.683
R586 VGND.n269 VGND.n268 462.683
R587 VGND.n268 VGND.n267 462.683
R588 VGND.n259 VGND.n40 462.683
R589 VGND.n261 VGND.n259 462.683
R590 VGND.n183 VGND.n182 411.555
R591 VGND.n180 VGND.n73 294.776
R592 VGND.n99 VGND.n98 294.776
R593 VGND.n130 VGND.n129 294.776
R594 VGND.n289 VGND.n20 294.776
R595 VGND.n212 VGND.n211 292.5
R596 VGND.n209 VGND.n187 292.5
R597 VGND.n209 VGND.n51 292.5
R598 VGND.n208 VGND.n207 292.5
R599 VGND.n206 VGND.n205 292.5
R600 VGND.n204 VGND.n203 292.5
R601 VGND.n55 VGND.n53 292.5
R602 VGND.n161 VGND.n78 280.32
R603 VGND.n300 VGND.n5 280.32
R604 VGND.n137 VGND.n77 268.425
R605 VGND.n145 VGND.n86 268.425
R606 VGND.n158 VGND.n157 268.425
R607 VGND.n121 VGND.n4 268.425
R608 VGND.n109 VGND.n104 268.425
R609 VGND.n108 VGND.n18 268.425
R610 VGND.n139 VGND.n137 268.274
R611 VGND.n123 VGND.n121 268.274
R612 VGND.n255 VGND.t7 266.909
R613 VGND.n145 VGND.n144 256.377
R614 VGND.n158 VGND.n86 256.377
R615 VGND.n128 VGND.n104 256.377
R616 VGND.n109 VGND.n108 256.377
R617 VGND.n162 VGND.n161 256
R618 VGND.n301 VGND.n300 256
R619 VGND.n48 VGND.n26 218.868
R620 VGND.n279 VGND.n1 211.994
R621 VGND.n208 VGND.n188 211.361
R622 VGND.n211 VGND.n210 211.361
R623 VGND.n205 VGND.n188 211.361
R624 VGND.n204 VGND.n196 211.137
R625 VGND.n196 VGND.n53 211.137
R626 VGND.n144 VGND.n98 209.695
R627 VGND.n157 VGND.n73 209.695
R628 VGND.n129 VGND.n128 209.695
R629 VGND.n20 VGND.n18 209.695
R630 VGND.t18 VGND.n70 202.168
R631 VGND.t24 VGND.n183 202.168
R632 VGND.n28 VGND.n1 199.947
R633 VGND.t0 VGND.n223 193.083
R634 VGND.n214 VGND.n213 156.988
R635 VGND.n226 VGND.n225 151.072
R636 VGND.n221 VGND.n220 146.25
R637 VGND.n219 VGND.n52 146.25
R638 VGND.n62 VGND.n61 146.25
R639 VGND.t22 VGND.t18 145.38
R640 VGND.t16 VGND.t22 145.38
R641 VGND.t16 VGND.t20 145.38
R642 VGND.t20 VGND.t24 145.38
R643 VGND.n278 VGND.n24 140.048
R644 VGND.n279 VGND.n278 135.906
R645 VGND.t39 VGND.n226 132.538
R646 VGND.n70 VGND.n51 130.614
R647 VGND.n222 VGND.n221 128.493
R648 VGND.n222 VGND.n52 128.493
R649 VGND.n28 VGND.n25 123.859
R650 VGND.n169 VGND.n62 119.719
R651 VGND.n219 VGND.n57 119.267
R652 VGND.n220 VGND.n54 119.267
R653 VGND.n61 VGND.n50 118.124
R654 VGND.n30 VGND.n29 117.475
R655 VGND.n234 VGND.n233 117.001
R656 VGND.n234 VGND.n49 117.001
R657 VGND.n242 VGND.n241 117.001
R658 VGND.n241 VGND.n49 117.001
R659 VGND.n246 VGND.n238 117.001
R660 VGND.n238 VGND.n49 117.001
R661 VGND.n29 VGND.n28 117.001
R662 VGND.n127 VGND.n126 117.001
R663 VGND.n126 VGND.n125 117.001
R664 VGND.n7 VGND.n5 117.001
R665 VGND.n9 VGND.n7 117.001
R666 VGND.n295 VGND.n294 117.001
R667 VGND.n294 VGND.n9 117.001
R668 VGND.n14 VGND.n13 117.001
R669 VGND.n13 VGND.n8 117.001
R670 VGND.n111 VGND.n110 117.001
R671 VGND.n111 VGND.n8 117.001
R672 VGND.n289 VGND.n19 117.001
R673 VGND.n282 VGND.n19 117.001
R674 VGND.n131 VGND.n130 117.001
R675 VGND.n132 VGND.n131 117.001
R676 VGND.n124 VGND.n123 117.001
R677 VGND.n125 VGND.n124 117.001
R678 VGND.n143 VGND.n142 117.001
R679 VGND.n142 VGND.n95 117.001
R680 VGND.n156 VGND.n155 117.001
R681 VGND.n155 VGND.n82 117.001
R682 VGND.n181 VGND.n180 117.001
R683 VGND.n182 VGND.n181 117.001
R684 VGND.n150 VGND.n149 117.001
R685 VGND.n149 VGND.n81 117.001
R686 VGND.n93 VGND.n87 117.001
R687 VGND.n93 VGND.n81 117.001
R688 VGND.n80 VGND.n78 117.001
R689 VGND.n82 VGND.n80 117.001
R690 VGND.n139 VGND.n138 117.001
R691 VGND.n138 VGND.n95 117.001
R692 VGND.n100 VGND.n99 117.001
R693 VGND.n133 VGND.n100 117.001
R694 VGND.n239 VGND.n227 117.001
R695 VGND.n254 VGND.n227 117.001
R696 VGND.n231 VGND.n224 117.001
R697 VGND.n254 VGND.n224 117.001
R698 VGND.n253 VGND.n252 117.001
R699 VGND.n254 VGND.n253 117.001
R700 VGND.n42 VGND.n37 117.001
R701 VGND.n274 VGND.n37 117.001
R702 VGND.n266 VGND.n265 117.001
R703 VGND.n265 VGND.n264 117.001
R704 VGND.n257 VGND.n44 117.001
R705 VGND.n264 VGND.n257 117.001
R706 VGND.n270 VGND.n35 117.001
R707 VGND.n274 VGND.n35 117.001
R708 VGND.n263 VGND.n262 117.001
R709 VGND.n264 VGND.n263 117.001
R710 VGND.n24 VGND.n21 117.001
R711 VGND.n281 VGND.n21 117.001
R712 VGND.n273 VGND.n272 117.001
R713 VGND.n274 VGND.n273 117.001
R714 VGND.n260 VGND.n26 117.001
R715 VGND.n280 VGND.n279 117.001
R716 VGND.n281 VGND.n280 117.001
R717 VGND.n218 VGND.n217 110.727
R718 VGND.n218 VGND.n62 101.944
R719 VGND.n262 VGND.n261 89.224
R720 VGND.n262 VGND.n45 89.224
R721 VGND.n243 VGND.n239 89.224
R722 VGND.n242 VGND.n232 89.224
R723 VGND.n245 VGND.n242 89.224
R724 VGND.n246 VGND.n245 89.224
R725 VGND.n252 VGND.n251 89.224
R726 VGND.n251 VGND.n231 89.224
R727 VGND.n243 VGND.n231 89.224
R728 VGND.n233 VGND.n232 89.224
R729 VGND.n267 VGND.n44 89.224
R730 VGND.n271 VGND.n270 89.224
R731 VGND.n270 VGND.n269 89.224
R732 VGND.n269 VGND.n42 89.224
R733 VGND.n266 VGND.n45 89.224
R734 VGND.n267 VGND.n266 89.224
R735 VGND.n40 VGND.n24 89.224
R736 VGND.n272 VGND.n40 89.224
R737 VGND.n272 VGND.n271 89.224
R738 VGND.n261 VGND.n260 89.224
R739 VGND.n64 VGND.t48 85.9987
R740 VGND.n151 VGND.n87 85.0829
R741 VGND.n87 VGND.n77 85.0829
R742 VGND.n157 VGND.n156 85.0829
R743 VGND.n150 VGND.n86 85.0829
R744 VGND.n144 VGND.n143 85.0829
R745 VGND.n14 VGND.n4 85.0829
R746 VGND.n15 VGND.n14 85.0829
R747 VGND.n110 VGND.n109 85.0829
R748 VGND.n295 VGND.n18 85.0829
R749 VGND.n128 VGND.n127 85.0829
R750 VGND.n168 VGND.t47 85.0821
R751 VGND.n136 VGND.n99 84.9588
R752 VGND.n130 VGND.n103 84.9588
R753 VGND.n180 VGND.n179 84.6953
R754 VGND.n290 VGND.n289 84.6953
R755 VGND.n185 VGND.t4 84.1654
R756 VGND.n189 VGND.t2 84.1654
R757 VGND.n191 VGND.t1 84.1654
R758 VGND.n193 VGND.t3 84.1654
R759 VGND.n197 VGND.t46 84.1654
R760 VGND.n201 VGND.t45 84.1654
R761 VGND.n199 VGND.t15 84.1654
R762 VGND.t34 VGND.n8 83.677
R763 VGND.t9 VGND.n9 83.677
R764 VGND.n281 VGND.t43 83.677
R765 VGND.n125 VGND.t34 79.9216
R766 VGND.t9 VGND.n8 79.9216
R767 VGND.n151 VGND.n92 66.6518
R768 VGND.n118 VGND.n15 66.6518
R769 VGND.n132 VGND.t26 65.3691
R770 VGND.n125 VGND.t26 65.3691
R771 VGND.t11 VGND.n9 65.3691
R772 VGND.t11 VGND.n282 65.3691
R773 VGND.n153 VGND.n152 64.7759
R774 VGND.n297 VGND.n296 64.7759
R775 VGND.n152 VGND.n151 63.1207
R776 VGND.n297 VGND.n15 63.1207
R777 VGND.n141 VGND.n92 61.2449
R778 VGND.n118 VGND.n105 61.2449
R779 VGND.n278 VGND.n277 60.6431
R780 VGND.t33 VGND.t43 60.5574
R781 VGND.n156 VGND.n153 58.5793
R782 VGND.n143 VGND.n141 58.5793
R783 VGND.n296 VGND.n295 58.5793
R784 VGND.n127 VGND.n105 58.5793
R785 VGND.n217 VGND.n216 58.5005
R786 VGND.n216 VGND.t16 58.5005
R787 VGND.n215 VGND.n214 58.5005
R788 VGND.t16 VGND.n215 58.5005
R789 VGND.n151 VGND.n150 54.2123
R790 VGND.n110 VGND.n15 54.2123
R791 VGND.n277 VGND.n276 54.1382
R792 VGND.n282 VGND.n281 47.0612
R793 VGND.n291 VGND.n290 41.7862
R794 VGND.t11 VGND.n291 41.7862
R795 VGND.n292 VGND.n20 41.7862
R796 VGND.n292 VGND.t11 41.7862
R797 VGND.n129 VGND.n102 41.7862
R798 VGND.n102 VGND.t26 41.7862
R799 VGND.n103 VGND.n101 41.7862
R800 VGND.n101 VGND.t26 41.7862
R801 VGND.n179 VGND.n72 41.7862
R802 VGND.n72 VGND.t37 41.7862
R803 VGND.n136 VGND.n135 41.7862
R804 VGND.n135 VGND.t31 41.7862
R805 VGND.n134 VGND.n98 41.7862
R806 VGND.t31 VGND.n134 41.7862
R807 VGND.n73 VGND.n71 41.7862
R808 VGND.n71 VGND.t37 41.7862
R809 VGND.n196 VGND.n51 40.6828
R810 VGND.n210 VGND.n51 40.571
R811 VGND.n188 VGND.n51 40.571
R812 VGND.n119 VGND.n118 34.4123
R813 VGND.t34 VGND.n119 34.4123
R814 VGND.n298 VGND.n297 34.4123
R815 VGND.t9 VGND.n298 34.4123
R816 VGND.n108 VGND.n10 34.4123
R817 VGND.t9 VGND.n10 34.4123
R818 VGND.n113 VGND.n104 34.4123
R819 VGND.t34 VGND.n113 34.4123
R820 VGND.n121 VGND.n120 34.4123
R821 VGND.n120 VGND.t34 34.4123
R822 VGND.n300 VGND.n299 34.4123
R823 VGND.n299 VGND.t9 34.4123
R824 VGND.n147 VGND.n92 34.4123
R825 VGND.n147 VGND.t28 34.4123
R826 VGND.n152 VGND.n83 34.4123
R827 VGND.t5 VGND.n83 34.4123
R828 VGND.n161 VGND.n160 34.4123
R829 VGND.n160 VGND.t5 34.4123
R830 VGND.n137 VGND.n96 34.4123
R831 VGND.t28 VGND.n96 34.4123
R832 VGND.n146 VGND.n145 34.4123
R833 VGND.t28 VGND.n146 34.4123
R834 VGND.n159 VGND.n158 34.4123
R835 VGND.t5 VGND.n159 34.4123
R836 VGND.n277 VGND.n23 34.4123
R837 VGND.n23 VGND.t43 34.4123
R838 VGND.n22 VGND.n1 34.4123
R839 VGND.n22 VGND.t43 34.4123
R840 VGND.n220 VGND.n219 32.0858
R841 VGND.n225 VGND.n34 30.9573
R842 VGND.n220 VGND.n55 28.5224
R843 VGND.n212 VGND.n187 22.5938
R844 VGND.n207 VGND.n187 22.5938
R845 VGND.n207 VGND.n206 22.5938
R846 VGND.n203 VGND.n55 22.5079
R847 VGND.n48 VGND.n30 21.964
R848 VGND.n136 VGND.t32 21.1687
R849 VGND.n179 VGND.t38 21.1687
R850 VGND.n103 VGND.t27 21.1687
R851 VGND.n290 VGND.t12 21.1687
R852 VGND.n213 VGND.n212 19.8448
R853 VGND.n223 VGND.n50 18.7528
R854 VGND.t33 VGND.n30 18.4903
R855 VGND.n153 VGND.n74 18.297
R856 VGND.n141 VGND.n140 18.297
R857 VGND.n296 VGND.n17 18.297
R858 VGND.n122 VGND.n105 18.297
R859 VGND.n69 VGND.n67 18.2817
R860 VGND.n183 VGND.n69 18.2817
R861 VGND.n195 VGND.n68 18.2817
R862 VGND.n70 VGND.n68 18.2817
R863 VGND.n57 VGND.t42 17.4005
R864 VGND.n57 VGND.t14 17.4005
R865 VGND.n54 VGND.t8 17.4005
R866 VGND.n54 VGND.t49 17.4005
R867 VGND.n88 VGND.t30 17.3591
R868 VGND.n165 VGND.t36 17.3591
R869 VGND.n114 VGND.t50 17.3591
R870 VGND.n283 VGND.t13 17.3591
R871 VGND.n250 VGND.n249 17.2064
R872 VGND.n249 VGND.t39 17.2064
R873 VGND.n244 VGND.n237 17.2064
R874 VGND.t39 VGND.n237 17.2064
R875 VGND.n248 VGND.n247 17.2064
R876 VGND.t39 VGND.n248 17.2064
R877 VGND.n230 VGND.n228 17.2064
R878 VGND.n228 VGND.n34 17.2064
R879 VGND.n43 VGND.n27 17.2064
R880 VGND.t33 VGND.n27 17.2064
R881 VGND.n268 VGND.n31 17.2064
R882 VGND.t33 VGND.n31 17.2064
R883 VGND.n41 VGND.n32 17.2064
R884 VGND.t33 VGND.n32 17.2064
R885 VGND.n259 VGND.n33 17.2064
R886 VGND.t33 VGND.n33 17.2064
R887 VGND.n276 VGND.n275 17.2064
R888 VGND.n275 VGND.t33 17.2064
R889 VGND.n1 VGND.t44 16.6948
R890 VGND.n152 VGND.t6 16.6948
R891 VGND.n92 VGND.t29 16.6948
R892 VGND.n118 VGND.t35 16.6948
R893 VGND.n297 VGND.t10 16.6948
R894 VGND.n206 VGND.n195 11.7696
R895 VGND.n203 VGND.n195 10.8247
R896 VGND.n175 VGND.t25 10.6446
R897 VGND.n174 VGND.n172 8.96117
R898 VGND.n174 VGND.n173 8.90463
R899 VGND.n223 VGND.n222 8.88039
R900 VGND.n179 VGND.n74 8.08353
R901 VGND.n140 VGND.n136 8.08353
R902 VGND.n122 VGND.n103 8.08353
R903 VGND.n290 VGND.n17 8.08353
R904 VGND.n276 VGND.n25 6.50542
R905 VGND.n115 VGND 6.13208
R906 VGND.n219 VGND.n218 5.1205
R907 VGND.n185 VGND.n184 4.68598
R908 VGND.n170 VGND.n169 4.6505
R909 VGND.n212 VGND.n186 4.6505
R910 VGND.n190 VGND.n187 4.6505
R911 VGND.n207 VGND.n192 4.6505
R912 VGND.n206 VGND.n194 4.6505
R913 VGND.n203 VGND.n202 4.6505
R914 VGND.n200 VGND.n55 4.6505
R915 VGND.n3 VGND 3.83932
R916 VGND.n117 VGND.n16 3.27485
R917 VGND.n91 VGND.n75 3.27485
R918 VGND.n220 VGND.n56 3.1005
R919 VGND.n219 VGND.n60 3.1005
R920 VGND.n63 VGND.n62 3.1005
R921 VGND.n78 VGND.n74 3.08756
R922 VGND.n140 VGND.n139 3.08756
R923 VGND.n17 VGND.n5 3.08756
R924 VGND.n123 VGND.n122 3.08756
R925 VGND.n213 VGND.n184 2.74949
R926 VGND.n285 VGND 1.89195
R927 VGND.n2 VGND 1.81103
R928 VGND.n172 VGND.t19 1.7405
R929 VGND.n172 VGND.t23 1.7405
R930 VGND.n173 VGND.t17 1.7405
R931 VGND.n173 VGND.t21 1.7405
R932 VGND.n303 VGND.n1 1.64558
R933 VGND.n167 VGND.n75 1.55665
R934 VGND.n285 VGND.n16 1.55665
R935 VGND.n91 VGND.n90 1.43327
R936 VGND.n117 VGND.n116 1.43327
R937 VGND.t7 VGND.t0 1.13628
R938 VGND.n223 VGND.n51 1.13628
R939 VGND.n65 VGND.n64 1.02133
R940 VGND.n89 VGND 0.931775
R941 VGND.n217 VGND.n66 0.9305
R942 VGND.n284 VGND 0.893921
R943 VGND.n116 VGND 0.875052
R944 VGND.n179 VGND.n178 0.846996
R945 VGND.n290 VGND.n288 0.845955
R946 VGND.n168 VGND 0.705857
R947 VGND.n304 VGND.n303 0.698599
R948 VGND.n176 VGND 0.672517
R949 VGND.n152 VGND.n75 0.664786
R950 VGND.n92 VGND.n91 0.664786
R951 VGND.n297 VGND.n16 0.664786
R952 VGND.n118 VGND.n117 0.664786
R953 VGND.n76 VGND 0.659154
R954 VGND.n304 VGND 0.648552
R955 VGND.n164 VGND 0.584663
R956 VGND.n177 VGND.n171 0.576446
R957 VGND.n177 VGND.n176 0.563
R958 VGND.n90 VGND 0.55129
R959 VGND.n305 VGND.n304 0.448175
R960 VGND.n162 VGND.n77 0.376971
R961 VGND.n301 VGND.n4 0.376971
R962 VGND.n302 VGND.n2 0.372211
R963 VGND.n285 VGND.n284 0.342605
R964 VGND.n166 VGND 0.324058
R965 VGND.n283 VGND.n3 0.321553
R966 VGND.n284 VGND.n283 0.321553
R967 VGND.n115 VGND.n114 0.321553
R968 VGND.n114 VGND.n2 0.321553
R969 VGND.n302 VGND.n3 0.316289
R970 VGND.n198 VGND.n195 0.3105
R971 VGND VGND.n0 0.290066
R972 VGND.n116 VGND.n115 0.289974
R973 VGND.n167 VGND 0.286855
R974 VGND.n58 VGND 0.281364
R975 VGND.n305 VGND.n0 0.248454
R976 VGND VGND.n177 0.235626
R977 VGND.n59 VGND 0.207231
R978 VGND.n286 VGND 0.205536
R979 VGND VGND.n56 0.200274
R980 VGND.n171 VGND 0.15335
R981 VGND.n186 VGND 0.146412
R982 VGND.n190 VGND 0.145792
R983 VGND.n192 VGND 0.145792
R984 VGND.n194 VGND 0.145792
R985 VGND VGND.n200 0.144985
R986 VGND.n163 VGND.n162 0.133357
R987 VGND.n302 VGND.n301 0.133357
R988 VGND.n66 VGND.n65 0.128645
R989 VGND.n165 VGND.n164 0.120692
R990 VGND.n166 VGND.n165 0.120692
R991 VGND.n89 VGND.n88 0.120692
R992 VGND.n88 VGND.n76 0.120692
R993 VGND.n163 VGND.n0 0.111589
R994 VGND.n303 VGND.n302 0.111589
R995 VGND.n60 VGND.n59 0.104667
R996 VGND.n202 VGND.n198 0.099378
R997 VGND VGND.n56 0.0954074
R998 VGND.n59 VGND.n58 0.0854359
R999 VGND.n178 VGND.n167 0.081623
R1000 VGND.n178 VGND 0.081623
R1001 VGND.n65 VGND 0.066858
R1002 VGND.n288 VGND.n287 0.063
R1003 VGND.n288 VGND.n286 0.0626302
R1004 VGND.n175 VGND.n174 0.0610124
R1005 VGND.n287 VGND 0.0540072
R1006 VGND.n286 VGND.n285 0.0540072
R1007 VGND.n163 VGND.n76 0.0537869
R1008 VGND.n167 VGND.n166 0.0493048
R1009 VGND.n198 VGND 0.0469135
R1010 VGND.n171 VGND.n66 0.0463595
R1011 VGND.n164 VGND.n163 0.0453207
R1012 VGND.n287 VGND 0.0445089
R1013 VGND.n90 VGND.n89 0.0413367
R1014 VGND.n189 VGND.n186 0.0346615
R1015 VGND.n191 VGND.n190 0.0346615
R1016 VGND.n193 VGND.n192 0.0346615
R1017 VGND.n197 VGND.n194 0.0346615
R1018 VGND.n202 VGND.n201 0.0346615
R1019 VGND.n200 VGND.n199 0.0346615
R1020 VGND.n65 VGND.n60 0.0290494
R1021 VGND VGND.n185 0.0287258
R1022 VGND VGND.n189 0.0276739
R1023 VGND VGND.n191 0.0276739
R1024 VGND VGND.n193 0.0276739
R1025 VGND VGND.n197 0.0276739
R1026 VGND.n201 VGND 0.0276739
R1027 VGND.n199 VGND 0.0276739
R1028 VGND VGND.n305 0.024
R1029 VGND.n176 VGND.n175 0.0239099
R1030 VGND.n170 VGND.n168 0.0190048
R1031 VGND.n65 VGND 0.0120304
R1032 VGND.n58 VGND 0.00975926
R1033 VGND.n64 VGND.n63 0.00495493
R1034 VGND.n63 VGND 0.00495493
R1035 VGND VGND.n170 0.00417012
R1036 ua[0].n2 ua[0].t2 899.324
R1037 ua[0].n3 ua[0].t2 898.659
R1038 ua[0].t1 ua[0].n2 898.442
R1039 ua[0].n3 ua[0].t1 897.754
R1040 ua[0].n0 ua[0].t0 895.625
R1041 ua[0].n0 ua[0].t3 894.172
R1042 ua[0].n1 ua[0].n0 6.30807
R1043 ua[0].n2 ua[0].n1 5.39021
R1044 ua[0].n4 ua[0].n3 5.38653
R1045 ua[0].n4 ua[0].n1 5.11108
R1046 ua[0] ua[0].n4 0.870692
R1047 X_TIMER.X_COMP_P_TOP.tail.n0 X_TIMER.X_COMP_P_TOP.tail.t5 28.3038
R1048 X_TIMER.X_COMP_P_TOP.tail.n2 X_TIMER.X_COMP_P_TOP.tail.t0 28.2925
R1049 X_TIMER.X_COMP_P_TOP.tail.n0 X_TIMER.X_COMP_P_TOP.tail.t3 28.0955
R1050 X_TIMER.X_COMP_P_TOP.tail.n1 X_TIMER.X_COMP_P_TOP.tail.t6 28.0955
R1051 X_TIMER.X_COMP_P_TOP.tail.n1 X_TIMER.X_COMP_P_TOP.tail.t1 28.0955
R1052 X_TIMER.X_COMP_P_TOP.tail.n3 X_TIMER.X_COMP_P_TOP.tail.t7 28.0921
R1053 X_TIMER.X_COMP_P_TOP.tail.n3 X_TIMER.X_COMP_P_TOP.tail.t2 28.0842
R1054 X_TIMER.X_COMP_P_TOP.tail.n2 X_TIMER.X_COMP_P_TOP.tail.t8 28.0724
R1055 X_TIMER.X_COMP_P_TOP.tail X_TIMER.X_COMP_P_TOP.tail.t4 23.519
R1056 X_TIMER.X_COMP_P_TOP.tail.n3 X_TIMER.X_COMP_P_TOP.tail.n2 0.417167
R1057 X_TIMER.X_COMP_P_TOP.tail.n1 X_TIMER.X_COMP_P_TOP.tail.n0 0.417167
R1058 X_TIMER.X_COMP_P_TOP.tail X_TIMER.X_COMP_P_TOP.tail.n3 0.387596
R1059 X_TIMER.X_COMP_P_TOP.tail X_TIMER.X_COMP_P_TOP.tail.n1 0.384638
R1060 X_TIMER.X_COMP_P_TOP.latch_right.n2 X_TIMER.X_COMP_P_TOP.latch_right.t7 114.778
R1061 X_TIMER.X_COMP_P_TOP.latch_right.n2 X_TIMER.X_COMP_P_TOP.latch_right.t8 106.572
R1062 X_TIMER.X_COMP_P_TOP.latch_right.n3 X_TIMER.X_COMP_P_TOP.latch_right.t3 28.4736
R1063 X_TIMER.X_COMP_P_TOP.latch_right.n3 X_TIMER.X_COMP_P_TOP.latch_right.t6 28.057
R1064 X_TIMER.X_COMP_P_TOP.latch_right.n4 X_TIMER.X_COMP_P_TOP.latch_right.t5 27.8467
R1065 X_TIMER.X_COMP_P_TOP.latch_right.n4 X_TIMER.X_COMP_P_TOP.latch_right.t4 27.4301
R1066 X_TIMER.X_COMP_P_TOP.latch_right.n0 X_TIMER.X_COMP_P_TOP.latch_right.t2 22.0141
R1067 X_TIMER.X_COMP_P_TOP.latch_right.n5 X_TIMER.X_COMP_P_TOP.latch_right.t0 20.4334
R1068 X_TIMER.X_COMP_P_TOP.latch_right.n6 X_TIMER.X_COMP_P_TOP.latch_right.n5 13.8274
R1069 X_TIMER.X_COMP_P_TOP.latch_right.n1 X_TIMER.X_COMP_P_TOP.latch_right.n0 0.582966
R1070 X_TIMER.X_COMP_P_TOP.latch_right.n1 X_TIMER.X_COMP_P_TOP.latch_right.n2 1.69623
R1071 X_TIMER.X_COMP_P_TOP.latch_right.n1 X_TIMER.X_COMP_P_TOP.latch_right.t1 95.1763
R1072 X_TIMER.X_COMP_P_TOP.latch_right X_TIMER.X_COMP_P_TOP.latch_right.n0 0.612947
R1073 X_TIMER.X_COMP_P_TOP.latch_right.n6 X_TIMER.X_COMP_P_TOP.latch_right.n3 0.418903
R1074 X_TIMER.X_COMP_P_TOP.latch_right.n5 X_TIMER.X_COMP_P_TOP.latch_right.n4 0.210569
R1075 X_TIMER.X_COMP_P_TOP.latch_right X_TIMER.X_COMP_P_TOP.latch_right.n6 0.0977222
R1076 X_TIMER.X_COMP_P_BOTTOM.tail.n3 X_TIMER.X_COMP_P_BOTTOM.tail.t2 28.3038
R1077 X_TIMER.X_COMP_P_BOTTOM.tail.n0 X_TIMER.X_COMP_P_BOTTOM.tail.t6 28.2925
R1078 X_TIMER.X_COMP_P_BOTTOM.tail.n5 X_TIMER.X_COMP_P_BOTTOM.tail.t5 28.0955
R1079 X_TIMER.X_COMP_P_BOTTOM.tail.n4 X_TIMER.X_COMP_P_BOTTOM.tail.t0 28.0955
R1080 X_TIMER.X_COMP_P_BOTTOM.tail.n3 X_TIMER.X_COMP_P_BOTTOM.tail.t4 28.0955
R1081 X_TIMER.X_COMP_P_BOTTOM.tail.n2 X_TIMER.X_COMP_P_BOTTOM.tail.t1 28.0921
R1082 X_TIMER.X_COMP_P_BOTTOM.tail.n1 X_TIMER.X_COMP_P_BOTTOM.tail.t7 28.0842
R1083 X_TIMER.X_COMP_P_BOTTOM.tail.n0 X_TIMER.X_COMP_P_BOTTOM.tail.t3 28.0724
R1084 X_TIMER.X_COMP_P_BOTTOM.tail X_TIMER.X_COMP_P_BOTTOM.tail.t8 23.519
R1085 X_TIMER.X_COMP_P_BOTTOM.tail X_TIMER.X_COMP_P_BOTTOM.tail.n2 0.387596
R1086 X_TIMER.X_COMP_P_BOTTOM.tail X_TIMER.X_COMP_P_BOTTOM.tail.n5 0.384638
R1087 X_TIMER.X_COMP_P_BOTTOM.tail.n5 X_TIMER.X_COMP_P_BOTTOM.tail.n4 0.208833
R1088 X_TIMER.X_COMP_P_BOTTOM.tail.n4 X_TIMER.X_COMP_P_BOTTOM.tail.n3 0.208833
R1089 X_TIMER.X_COMP_P_BOTTOM.tail.n2 X_TIMER.X_COMP_P_BOTTOM.tail.n1 0.208833
R1090 X_TIMER.X_COMP_P_BOTTOM.tail.n1 X_TIMER.X_COMP_P_BOTTOM.tail.n0 0.208833
R1091 X_TIMER.X_SR_LATCH.IN_S.n0 X_TIMER.X_SR_LATCH.IN_S.t3 565.548
R1092 X_TIMER.X_SR_LATCH.IN_S.n0 X_TIMER.X_SR_LATCH.IN_S.t2 250.073
R1093 X_TIMER.X_SR_LATCH.IN_S X_TIMER.X_SR_LATCH.IN_S.n0 161.315
R1094 X_TIMER.X_SR_LATCH.IN_S X_TIMER.X_SR_LATCH.IN_S.t0 32.8039
R1095 X_TIMER.X_SR_LATCH.IN_S.n2 X_TIMER.X_SR_LATCH.IN_S.n1 18.3183
R1096 X_TIMER.X_SR_LATCH.IN_S.n2 X_TIMER.X_SR_LATCH.IN_S.t1 17.6591
R1097 X_TIMER.X_SR_LATCH.IN_S X_TIMER.X_SR_LATCH.IN_S.n2 10.7227
R1098 X_TIMER.X_SR_LATCH.IN_S.n1 X_TIMER.X_SR_LATCH.IN_S 5.53461
R1099 X_TIMER.X_SR_LATCH.IN_S.n1 X_TIMER.X_SR_LATCH.IN_S 3.78946
R1100 X_TIMER.X_COMP_P_TOP.out_left.n1 X_TIMER.X_COMP_P_TOP.out_left.t3 146.125
R1101 X_TIMER.X_COMP_P_TOP.out_left.n0 X_TIMER.X_COMP_P_TOP.out_left.t1 29.4286
R1102 X_TIMER.X_COMP_P_TOP.out_left X_TIMER.X_COMP_P_TOP.out_left.t2 20.2226
R1103 X_TIMER.X_COMP_P_TOP.out_left X_TIMER.X_COMP_P_TOP.out_left.n0 11.6041
R1104 X_TIMER.X_COMP_P_TOP.out_left.n0 X_TIMER.X_COMP_P_TOP.out_left.n1 1.08492
R1105 X_TIMER.X_COMP_P_TOP.out_left.t0 X_TIMER.X_COMP_P_TOP.out_left.n1 144.458
R1106 X_TIMER.X_SR_LATCH.inv_0.vin X_TIMER.X_SR_LATCH.IN_R.t3 411.07
R1107 X_TIMER.X_SR_LATCH.inv_0.vin X_TIMER.X_SR_LATCH.IN_R.t2 400.375
R1108 X_TIMER.X_SR_LATCH.IN_R.n0 X_TIMER.X_SR_LATCH.inv_0.vin 34.7689
R1109 X_TIMER.X_COMP_P_TOP.vout X_TIMER.X_SR_LATCH.IN_R.t0 32.8039
R1110 X_TIMER.X_SR_LATCH.IN_R.n0 X_TIMER.X_SR_LATCH.IN_R.t1 21.6505
R1111 X_TIMER.X_COMP_P_TOP.vout X_TIMER.X_SR_LATCH.IN_R.n0 6.73127
R1112 ui_in[0].n0 ui_in[0].t0 565.548
R1113 ui_in[0].n0 ui_in[0].t1 250.073
R1114 ui_in[0].n2 ui_in[0].n0 161.855
R1115 ui_in[0] ui_in[0].n2 6.27244
R1116 ui_in[0].n1 ui_in[0] 0.163962
R1117 ui_in[0].n2 ui_in[0].n1 0.0838333
R1118 ui_in[0].n1 ui_in[0] 0.0305926
R1119 ua[1].t1 ua[1].n1 899.351
R1120 ua[1].n2 ua[1].t1 898.639
R1121 ua[1].t0 ua[1].n1 898.442
R1122 ua[1].n2 ua[1].t0 897.758
R1123 ua[1].n0 ua[1].t3 894.928
R1124 ua[1].n0 ua[1].t2 893.475
R1125 ua[1].n3 ua[1].n1 10.0477
R1126 ua[1].n4 ua[1].n3 5.65194
R1127 ua[1].n3 ua[1].n2 4.91594
R1128 ua[1].n4 ua[1].n0 1.38866
R1129 ua[1] ua[1].n4 0.680788
R1130 X_TIMER.X_COMP_P_BOTTOM.latch_left.n1 X_TIMER.X_COMP_P_BOTTOM.latch_left.t7 114.778
R1131 X_TIMER.X_COMP_P_BOTTOM.latch_left.n1 X_TIMER.X_COMP_P_BOTTOM.latch_left.t8 106.572
R1132 X_TIMER.X_COMP_P_BOTTOM.latch_left.n2 X_TIMER.X_COMP_P_BOTTOM.latch_left.t1 95.1712
R1133 X_TIMER.X_COMP_P_BOTTOM.latch_left.n0 X_TIMER.X_COMP_P_BOTTOM.latch_left.t3 28.4943
R1134 X_TIMER.X_COMP_P_BOTTOM.latch_left.n0 X_TIMER.X_COMP_P_BOTTOM.latch_left.t4 28.0776
R1135 X_TIMER.X_COMP_P_BOTTOM.latch_left.n4 X_TIMER.X_COMP_P_BOTTOM.latch_left.t5 27.8805
R1136 X_TIMER.X_COMP_P_BOTTOM.latch_left.n4 X_TIMER.X_COMP_P_BOTTOM.latch_left.t6 27.4638
R1137 X_TIMER.X_COMP_P_BOTTOM.latch_left.n3 X_TIMER.X_COMP_P_BOTTOM.latch_left.t2 22.0141
R1138 X_TIMER.X_COMP_P_BOTTOM.latch_left.n5 X_TIMER.X_COMP_P_BOTTOM.latch_left.t0 20.6741
R1139 X_TIMER.X_COMP_P_BOTTOM.latch_left.n6 X_TIMER.X_COMP_P_BOTTOM.latch_left.n5 13.8226
R1140 X_TIMER.X_COMP_P_BOTTOM.latch_left.n2 X_TIMER.X_COMP_P_BOTTOM.latch_left.n1 1.72733
R1141 X_TIMER.X_COMP_P_BOTTOM.latch_left.n6 X_TIMER.X_COMP_P_BOTTOM.latch_left.n3 0.632444
R1142 X_TIMER.X_COMP_P_BOTTOM.latch_left.n3 X_TIMER.X_COMP_P_BOTTOM.latch_left.n2 0.599169
R1143 X_TIMER.X_COMP_P_BOTTOM.latch_left X_TIMER.X_COMP_P_BOTTOM.latch_left.n0 0.403278
R1144 X_TIMER.X_COMP_P_BOTTOM.latch_left.n5 X_TIMER.X_COMP_P_BOTTOM.latch_left.n4 0.280014
R1145 X_TIMER.X_COMP_P_BOTTOM.latch_left X_TIMER.X_COMP_P_BOTTOM.latch_left.n6 0.0855694
R1146 X_TIMER.X_COMP_P_BOTTOM.out_left.n0 X_TIMER.X_COMP_P_BOTTOM.out_left.t1 29.4286
R1147 X_TIMER.X_COMP_P_BOTTOM.out_left X_TIMER.X_COMP_P_BOTTOM.out_left.t2 20.2226
R1148 X_TIMER.X_COMP_P_BOTTOM.out_left X_TIMER.X_COMP_P_BOTTOM.out_left.n0 11.6041
R1149 X_TIMER.X_COMP_P_BOTTOM.out_left.n0 X_TIMER.X_COMP_P_BOTTOM.out_left.n1 1.08492
R1150 X_TIMER.X_COMP_P_BOTTOM.out_left.t3 X_TIMER.X_COMP_P_BOTTOM.out_left.n1 146.125
R1151 X_TIMER.X_COMP_P_BOTTOM.out_left.t0 X_TIMER.X_COMP_P_BOTTOM.out_left.n1 144.458
R1152 X_TIMER.X_COMP_P_TOP.latch_left.n0 X_TIMER.X_COMP_P_TOP.latch_left.t7 114.778
R1153 X_TIMER.X_COMP_P_TOP.latch_left.n0 X_TIMER.X_COMP_P_TOP.latch_left.t8 106.572
R1154 X_TIMER.X_COMP_P_TOP.latch_left.n1 X_TIMER.X_COMP_P_TOP.latch_left.t4 95.1712
R1155 X_TIMER.X_COMP_P_TOP.latch_left.n6 X_TIMER.X_COMP_P_TOP.latch_left.t3 28.4943
R1156 X_TIMER.X_COMP_P_TOP.latch_left.n6 X_TIMER.X_COMP_P_TOP.latch_left.t1 28.0776
R1157 X_TIMER.X_COMP_P_TOP.latch_left.n3 X_TIMER.X_COMP_P_TOP.latch_left.t0 27.8805
R1158 X_TIMER.X_COMP_P_TOP.latch_left.n3 X_TIMER.X_COMP_P_TOP.latch_left.t2 27.4638
R1159 X_TIMER.X_COMP_P_TOP.latch_left.n2 X_TIMER.X_COMP_P_TOP.latch_left.t5 22.0141
R1160 X_TIMER.X_COMP_P_TOP.latch_left.n4 X_TIMER.X_COMP_P_TOP.latch_left.t6 20.6741
R1161 X_TIMER.X_COMP_P_TOP.latch_left.n5 X_TIMER.X_COMP_P_TOP.latch_left.n4 13.8226
R1162 X_TIMER.X_COMP_P_TOP.latch_left.n1 X_TIMER.X_COMP_P_TOP.latch_left.n0 1.72733
R1163 X_TIMER.X_COMP_P_TOP.latch_left.n5 X_TIMER.X_COMP_P_TOP.latch_left.n2 0.632444
R1164 X_TIMER.X_COMP_P_TOP.latch_left.n2 X_TIMER.X_COMP_P_TOP.latch_left.n1 0.599169
R1165 X_TIMER.X_COMP_P_TOP.latch_left X_TIMER.X_COMP_P_TOP.latch_left.n6 0.403278
R1166 X_TIMER.X_COMP_P_TOP.latch_left.n4 X_TIMER.X_COMP_P_TOP.latch_left.n3 0.280014
R1167 X_TIMER.X_COMP_P_TOP.latch_left X_TIMER.X_COMP_P_TOP.latch_left.n5 0.0855694
R1168 ua[2].n1 ua[2].t1 10.6631
R1169 ua[2].n1 ua[2].n0 8.86659
R1170 ua[2].n3 ua[2].n2 8.86659
R1171 ua[2].n4 ua[2] 7.67213
R1172 ua[2].n0 ua[2].t3 1.7405
R1173 ua[2].n0 ua[2].t0 1.7405
R1174 ua[2].n2 ua[2].t2 1.7405
R1175 ua[2].n2 ua[2].t4 1.7405
R1176 ua[2] ua[2].n3 0.160394
R1177 ua[2].n3 ua[2].n1 0.0570371
R1178 ua[2].n4 ua[2] 0.0537667
R1179 ua[2] ua[2].n4 0.0448889
C0 ui_in[0] X_TIMER.X_SR_LATCH.IN_S 0.172333f
C1 X_TIMER.X_COMP_P_BOTTOM.out_left X_TIMER.X_COMP_P_BOTTOM.tail 0.004812f
C2 X_TIMER.q_sr a_1723_2994# 0.161311f
C3 X_TIMER.X_COMP_P_BOTTOM.latch_right X_TIMER.X_COMP_P_BOTTOM.out_left 0.142667f
C4 ui_in[0] uio_in[5] 0.010273f
C5 X_TIMER.q_sr X_TIMER.out_inv1 0.324343f
C6 X_TIMER.X_COMP_P_TOP.latch_left X_TIMER.X_COMP_P_TOP.tail 8.829929f
C7 a_1723_2994# X_TIMER.X_SR_LATCH.IN_S 0.001116f
C8 ua[1] VPWR 3.56896f
C9 X_TIMER.out_inv1 X_TIMER.X_SR_LATCH.IN_S 0.046905f
C10 X_TIMER.bias_2 X_TIMER.bias_1 0.013902f
C11 uo_out[0] uio_oe[4] 0.013858f
C12 a_1347_2994# VPWR 0.183384f
C13 ua[2] X_TIMER.qb_sr 9.87e-19
C14 ua[1] X_TIMER.v1p2 1.12448f
C15 X_TIMER.X_COMP_P_BOTTOM.out_left X_TIMER.v0p6 0.233377f
C16 ui_in[6] ui_in[0] 0.010273f
C17 X_TIMER.X_COMP_P_TOP.latch_right X_TIMER.bias_p 0.001093f
C18 uio_in[4] uio_in[5] 0.023797f
C19 ui_in[0] uio_in[6] 0.010273f
C20 uo_out[3] uo_out[0] 0.013858f
C21 uio_in[3] uio_in[2] 0.023797f
C22 uo_out[0] uio_out[3] 0.013858f
C23 uo_out[0] ua[1] 0.347629f
C24 X_TIMER.v1p2 VPWR 3.82833f
C25 ua[1] X_TIMER.out_inv3 0.21732f
C26 uio_out[1] uio_out[0] 0.023797f
C27 X_TIMER.X_COMP_P_BOTTOM.tail X_TIMER.X_SR_LATCH.IN_S 0.010782f
C28 uio_oe[4] uio_oe[3] 0.023797f
C29 uio_out[1] uio_out[2] 0.023797f
C30 X_TIMER.X_COMP_P_BOTTOM.latch_right X_TIMER.X_SR_LATCH.IN_S 1.00897f
C31 uo_out[0] uio_oe[0] 0.013858f
C32 a_1347_2994# X_TIMER.out_inv3 1.51e-20
C33 ui_in[0] X_TIMER.bias_3 6e-19
C34 X_TIMER.bias_n ua[0] 0.252991f
C35 uo_out[0] VPWR 8.46475f
C36 a_1347_2994# X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B 5.92e-20
C37 X_TIMER.out_inv3 VPWR 1.74376f
C38 X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B VPWR 0.767973f
C39 uo_out[0] X_TIMER.v1p2 0.150366f
C40 ui_in[0] X_TIMER.X_SR_LATCH.nand_0.drain_mna 0.016193f
C41 uio_oe[5] uio_oe[6] 0.023797f
C42 ui_in[0] ui_in[3] 0.010273f
C43 ua[2] X_TIMER.out_inv1 5.71e-19
C44 ui_in[4] ui_in[3] 0.023797f
C45 X_TIMER.v1p2 X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B 1.51e-19
C46 X_TIMER.v0p6 X_TIMER.X_SR_LATCH.IN_S 0.038925f
C47 uo_out[2] uo_out[1] 0.023797f
C48 ua[1] X_TIMER.bias_p 0.189287f
C49 uo_out[0] uio_oe[2] 0.013858f
C50 X_TIMER.q_sr X_TIMER.X_SR_LATCH.nand_0.IN_A 0.004227f
C51 uo_out[4] uo_out[5] 0.023797f
C52 X_TIMER.X_COMP_P_BOTTOM.latch_left X_TIMER.X_COMP_P_BOTTOM.tail 8.82799f
C53 uo_out[0] X_TIMER.out_inv3 1.32372f
C54 X_TIMER.X_COMP_P_BOTTOM.latch_right X_TIMER.X_COMP_P_BOTTOM.latch_left 5.38251f
C55 uo_out[0] X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B 7.62e-19
C56 X_TIMER.X_SR_LATCH.nand_0.IN_A X_TIMER.X_SR_LATCH.IN_S 0.199334f
C57 X_TIMER.bias_p VPWR 12.319201f
C58 ui_in[0] X_TIMER.qb_sr 4.29e-20
C59 X_TIMER.out_inv3 X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B 1.61e-19
C60 X_TIMER.bias_n X_TIMER.bias_2 0.069293f
C61 uo_out[0] uo_out[6] 0.013858f
C62 X_TIMER.v1p2 X_TIMER.bias_p 0.361027f
C63 X_TIMER.X_COMP_P_BOTTOM.latch_right ua[2] 0.011181f
C64 uio_oe[3] uio_oe[2] 0.023797f
C65 ua[7] VPWR 0.010285f
C66 a_1723_2994# X_TIMER.qb_sr 0.006959f
C67 uo_out[0] uio_oe[3] 0.013858f
C68 X_TIMER.X_COMP_P_BOTTOM.latch_left X_TIMER.v0p6 0.504304f
C69 X_TIMER.out_inv1 X_TIMER.qb_sr 0.002285f
C70 X_TIMER.bias_2 X_TIMER.bias_3 0.013902f
C71 uo_out[0] X_TIMER.bias_p 3.21e-19
C72 X_TIMER.X_COMP_P_TOP.latch_left X_TIMER.X_COMP_P_TOP.latch_right 5.38251f
C73 ui_in[0] ui_in[4] 0.010273f
C74 uo_out[0] uio_in[7] 0.023797f
C75 ui_in[0] ui_in[1] 0.034283f
C76 uo_out[0] uo_out[7] 0.013858f
C77 ui_in[6] ui_in[7] 0.023797f
C78 X_TIMER.X_COMP_P_TOP.out_left ua[0] 0.244712f
C79 ua[1] X_TIMER.X_COMP_P_BOTTOM.out_left 0.389294f
C80 ui_in[0] uio_in[4] 0.010273f
C81 uo_out[7] uo_out[6] 0.023797f
C82 X_TIMER.X_COMP_P_TOP.out_left X_TIMER.X_COMP_P_TOP.tail 0.006519f
C83 X_TIMER.X_COMP_P_BOTTOM.out_left VPWR 6.37052f
C84 ua[6] ua[2] 0.0564f
C85 X_TIMER.X_SR_LATCH.nand_0.IN_A X_TIMER.X_SR_LATCH.nand_0.drain_mna 0.001812f
C86 X_TIMER.X_COMP_P_TOP.latch_left ua[1] 0.071128f
C87 X_TIMER.bias_1 VPWR 0.387201f
C88 X_TIMER.v1p2 X_TIMER.X_COMP_P_BOTTOM.out_left 0.008724f
C89 X_TIMER.X_COMP_P_TOP.out_left X_TIMER.X_COMP_P_BOTTOM.tail 3.1e-21
C90 uio_out[6] uio_out[5] 0.023797f
C91 uo_out[0] uo_out[1] 0.037655f
C92 ui_in[0] rst_n 0.02398f
C93 X_TIMER.X_COMP_P_TOP.tail ua[0] 2.92045f
C94 uo_out[0] X_TIMER.X_COMP_P_BOTTOM.out_left 0.13262f
C95 X_TIMER.X_COMP_P_TOP.latch_left VPWR 1.81653f
C96 X_TIMER.out_inv3 X_TIMER.X_COMP_P_BOTTOM.out_left 0.013941f
C97 X_TIMER.q_sr a_1347_2994# 0.015256f
C98 ua[1] X_TIMER.X_SR_LATCH.IN_S 0.145485f
C99 uo_out[0] X_TIMER.bias_1 4.12e-19
C100 X_TIMER.X_COMP_P_TOP.latch_left X_TIMER.v1p2 1.33915f
C101 X_TIMER.X_SR_LATCH.nand_0.IN_A X_TIMER.qb_sr 3.76e-20
C102 uio_in[2] uio_in[1] 0.023797f
C103 X_TIMER.q_sr VPWR 0.845552f
C104 a_1347_2994# X_TIMER.X_SR_LATCH.IN_S 0.009427f
C105 ua[2] ua[3] 0.0564f
C106 X_TIMER.X_COMP_P_TOP.out_left X_TIMER.v0p6 6.4e-22
C107 X_TIMER.bias_2 ua[0] 0.248813f
C108 uio_out[2] uio_out[3] 0.023797f
C109 X_TIMER.q_sr X_TIMER.v1p2 7.67e-21
C110 ui_in[0] uio_in[0] 0.010273f
C111 VPWR X_TIMER.X_SR_LATCH.IN_S 3.47783f
C112 uo_out[3] uo_out[4] 0.023797f
C113 X_TIMER.v1p2 X_TIMER.X_SR_LATCH.IN_S 1.61e-19
C114 X_TIMER.X_COMP_P_BOTTOM.out_left X_TIMER.bias_p 0.793062f
C115 ui_in[0] X_TIMER.X_SR_LATCH.nand_0.IN_A 0.281221f
C116 uo_out[0] X_TIMER.q_sr 7.86e-20
C117 X_TIMER.q_sr X_TIMER.out_inv3 2.38e-20
C118 ui_in[7] ui_in[0] 0.010273f
C119 X_TIMER.bias_1 X_TIMER.bias_p 0.056605f
C120 ua[1] X_TIMER.X_COMP_P_BOTTOM.latch_left 1.35459f
C121 X_TIMER.bias_n ua[1] 0.065657f
C122 X_TIMER.X_COMP_P_BOTTOM.latch_right X_TIMER.X_COMP_P_BOTTOM.tail 8.89308f
C123 X_TIMER.q_sr X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B 0.313825f
C124 uo_out[0] X_TIMER.X_SR_LATCH.IN_S 0.110526f
C125 X_TIMER.out_inv3 X_TIMER.X_SR_LATCH.IN_S 0.177402f
C126 ui_in[0] uio_in[3] 0.010273f
C127 ua[5] ua[2] 0.0564f
C128 X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B X_TIMER.X_SR_LATCH.IN_S 0.476501f
C129 X_TIMER.X_SR_LATCH.nand_0.IN_A X_TIMER.out_inv1 1.05e-20
C130 ua[1] ua[2] 4.93575f
C131 X_TIMER.X_COMP_P_TOP.latch_left X_TIMER.bias_p 0.001028f
C132 X_TIMER.X_COMP_P_BOTTOM.latch_left VPWR 1.83951f
C133 X_TIMER.bias_n VPWR 0.014926f
C134 uo_out[0] uio_out[0] 0.013858f
C135 uo_out[0] uio_out[2] 0.013858f
C136 X_TIMER.v0p6 X_TIMER.X_COMP_P_BOTTOM.tail 2.67476f
C137 uo_out[0] uo_out[4] 0.013858f
C138 X_TIMER.X_COMP_P_BOTTOM.latch_right X_TIMER.v0p6 0.512754f
C139 clk ena 0.023797f
C140 uo_out[0] uio_oe[6] 0.013858f
C141 ua[2] VPWR 0.034427f
C142 uio_in[4] uio_in[3] 0.023797f
C143 VPWR X_TIMER.bias_3 0.050264f
C144 X_TIMER.X_COMP_P_TOP.out_left X_TIMER.X_COMP_P_TOP.latch_right 0.143103f
C145 X_TIMER.bias_p X_TIMER.X_SR_LATCH.IN_S 0.094554f
C146 uo_out[0] uio_out[6] 0.013858f
C147 uo_out[0] X_TIMER.X_COMP_P_BOTTOM.latch_left 2.39e-19
C148 X_TIMER.X_COMP_P_BOTTOM.latch_left X_TIMER.out_inv3 0.029394f
C149 X_TIMER.X_SR_LATCH.nand_0.drain_mna VPWR 0.006259f
C150 clk rst_n 0.023797f
C151 uio_out[7] uio_oe[0] 0.023797f
C152 uo_out[0] ua[2] 8.56e-19
C153 X_TIMER.X_COMP_P_TOP.latch_right ua[0] 0.515831f
C154 uo_out[0] X_TIMER.bias_3 4.12e-19
C155 X_TIMER.out_inv3 ua[2] 0.802431f
C156 ua[2] X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B 0.001066f
C157 a_1347_2994# X_TIMER.qb_sr 0.150907f
C158 uio_out[0] uo_out[7] 0.023797f
C159 ua[2] ua[4] 0.0564f
C160 X_TIMER.X_COMP_P_TOP.tail X_TIMER.X_COMP_P_TOP.latch_right 8.89421f
C161 X_TIMER.X_COMP_P_BOTTOM.latch_left X_TIMER.bias_p 5.57e-19
C162 X_TIMER.qb_sr VPWR 0.532257f
C163 X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B X_TIMER.X_SR_LATCH.nand_0.drain_mna 0.080424f
C164 ui_in[7] uio_in[0] 0.023797f
C165 uio_out[7] uo_out[0] 0.013858f
C166 ua[1] X_TIMER.X_COMP_P_TOP.out_left 0.161037f
C167 X_TIMER.v1p2 X_TIMER.qb_sr 1.78e-19
C168 uio_in[6] uio_in[7] 0.023797f
C169 X_TIMER.bias_p X_TIMER.bias_3 6.09e-20
C170 X_TIMER.X_COMP_P_TOP.out_left VPWR 6.35315f
C171 uo_out[0] X_TIMER.qb_sr 8.53e-19
C172 X_TIMER.X_COMP_P_BOTTOM.out_left X_TIMER.X_SR_LATCH.IN_S 1.35688f
C173 ui_in[0] VPWR 1.12481f
C174 ua[1] ua[0] 10.7429f
C175 X_TIMER.out_inv3 X_TIMER.qb_sr 6.26e-19
C176 X_TIMER.X_COMP_P_TOP.out_left X_TIMER.v1p2 0.450222f
C177 X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B X_TIMER.qb_sr 0.448959f
C178 uio_oe[5] uio_oe[4] 0.023797f
C179 ui_in[3] ui_in[2] 0.023797f
C180 ui_in[0] X_TIMER.v1p2 5.91e-19
C181 a_1723_2994# VPWR 0.182866f
C182 ua[1] X_TIMER.X_COMP_P_TOP.tail 0.010057f
C183 ua[0] VPWR 5.19898f
C184 X_TIMER.out_inv1 VPWR 0.970352f
C185 uo_out[0] ui_in[0] 19.736f
C186 X_TIMER.v1p2 ua[0] 1.45006f
C187 X_TIMER.v1p2 X_TIMER.out_inv1 1.53e-20
C188 ui_in[0] X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B 0.114999f
C189 X_TIMER.X_COMP_P_TOP.tail VPWR 5.0999f
C190 ua[1] X_TIMER.X_COMP_P_BOTTOM.tail 0.83649f
C191 uio_oe[0] uio_oe[1] 0.023797f
C192 uio_out[5] uio_out[4] 0.023797f
C193 X_TIMER.q_sr X_TIMER.X_SR_LATCH.IN_S 0.306057f
C194 X_TIMER.X_COMP_P_BOTTOM.latch_left X_TIMER.X_COMP_P_BOTTOM.out_left 0.84597f
C195 ua[1] X_TIMER.X_COMP_P_BOTTOM.latch_right 3.57597f
C196 X_TIMER.v1p2 X_TIMER.X_COMP_P_TOP.tail 0.827015f
C197 uo_out[0] X_TIMER.out_inv1 0.678948f
C198 ua[1] X_TIMER.bias_2 0.086205f
C199 a_1723_2994# X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B 0.006917f
C200 X_TIMER.X_COMP_P_BOTTOM.tail VPWR 5.61759f
C201 X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B X_TIMER.out_inv1 0.001405f
C202 X_TIMER.X_COMP_P_BOTTOM.out_left ua[2] 0.005338f
C203 X_TIMER.X_COMP_P_BOTTOM.latch_right VPWR 1.695f
C204 ui_in[0] ui_in[2] 0.010273f
C205 X_TIMER.X_COMP_P_TOP.out_left X_TIMER.bias_p 0.845436f
C206 uo_out[0] uio_out[1] 0.013858f
C207 ui_in[0] X_TIMER.bias_p 3.36e-19
C208 ui_in[6] ui_in[5] 0.023797f
C209 uio_oe[1] uio_oe[2] 0.023797f
C210 X_TIMER.bias_2 VPWR 0.165891f
C211 ua[1] X_TIMER.v0p6 1.37952f
C212 X_TIMER.X_COMP_P_TOP.latch_left X_TIMER.bias_n 0.001099f
C213 ui_in[0] uio_in[1] 0.010273f
C214 uo_out[0] uio_oe[1] 0.013858f
C215 X_TIMER.bias_1 X_TIMER.bias_3 0.06887f
C216 ui_in[1] ui_in[2] 0.023797f
C217 uo_out[0] uio_oe[5] 0.013858f
C218 ui_in[0] uio_in[7] 0.010273f
C219 X_TIMER.bias_2 X_TIMER.v1p2 2.52e-19
C220 uo_out[0] X_TIMER.X_COMP_P_BOTTOM.tail 3.93e-19
C221 uo_out[0] X_TIMER.X_COMP_P_BOTTOM.latch_right 4.16e-19
C222 ua[0] X_TIMER.bias_p 0.099567f
C223 X_TIMER.v0p6 VPWR 5.94014f
C224 X_TIMER.X_COMP_P_BOTTOM.latch_right X_TIMER.out_inv3 0.003058f
C225 X_TIMER.X_COMP_P_BOTTOM.latch_left X_TIMER.X_SR_LATCH.IN_S 0.262546f
C226 uio_out[3] uio_out[4] 0.023797f
C227 uo_out[0] uo_out[5] 0.013858f
C228 X_TIMER.v1p2 X_TIMER.v0p6 0.171548f
C229 X_TIMER.q_sr ua[2] 7.94e-19
C230 uio_in[5] uio_in[6] 0.023797f
C231 X_TIMER.X_COMP_P_TOP.tail X_TIMER.bias_p 0.870817f
C232 ui_in[0] uio_in[2] 0.010273f
C233 X_TIMER.X_SR_LATCH.nand_0.IN_A VPWR 0.448244f
C234 ua[2] X_TIMER.X_SR_LATCH.IN_S 0.274914f
C235 uo_out[0] X_TIMER.v0p6 0.431659f
C236 uo_out[5] uo_out[6] 0.023797f
C237 X_TIMER.q_sr X_TIMER.X_SR_LATCH.nand_0.drain_mna 5.16e-21
C238 X_TIMER.out_inv3 X_TIMER.v0p6 0.002838f
C239 X_TIMER.X_COMP_P_BOTTOM.tail X_TIMER.bias_p 0.869796f
C240 uo_out[3] uo_out[2] 0.023797f
C241 X_TIMER.X_COMP_P_BOTTOM.latch_right X_TIMER.bias_p 7.91e-19
C242 X_TIMER.X_SR_LATCH.nand_0.drain_mna X_TIMER.X_SR_LATCH.IN_S 0.008133f
C243 uo_out[0] X_TIMER.X_SR_LATCH.nand_0.IN_A 4.72e-20
C244 X_TIMER.X_COMP_P_TOP.out_left X_TIMER.X_COMP_P_BOTTOM.out_left 0.016634f
C245 X_TIMER.bias_2 X_TIMER.bias_p 0.069262f
C246 ua[1] X_TIMER.X_COMP_P_TOP.latch_right 0.090139f
C247 uo_out[0] uio_out[4] 0.013858f
C248 X_TIMER.X_SR_LATCH.nand_0.IN_A X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B 0.239207f
C249 ui_in[0] X_TIMER.bias_1 6e-19
C250 X_TIMER.q_sr X_TIMER.qb_sr 0.385679f
C251 X_TIMER.X_COMP_P_BOTTOM.latch_left ua[2] 0.011758f
C252 X_TIMER.v0p6 X_TIMER.bias_p 0.030094f
C253 ua[0] X_TIMER.X_COMP_P_BOTTOM.out_left 1e-20
C254 X_TIMER.X_COMP_P_BOTTOM.out_left X_TIMER.out_inv1 1.75e-19
C255 X_TIMER.bias_n X_TIMER.bias_3 0.013902f
C256 X_TIMER.X_COMP_P_TOP.latch_right VPWR 1.65893f
C257 X_TIMER.qb_sr X_TIMER.X_SR_LATCH.IN_S 0.340841f
C258 X_TIMER.X_COMP_P_TOP.latch_left X_TIMER.X_COMP_P_TOP.out_left 0.846923f
C259 uio_in[0] uio_in[1] 0.023797f
C260 ui_in[0] ui_in[5] 0.010273f
C261 X_TIMER.v1p2 X_TIMER.X_COMP_P_TOP.latch_right 3.53509f
C262 X_TIMER.X_COMP_P_TOP.tail X_TIMER.X_COMP_P_BOTTOM.out_left 3.1e-21
C263 ui_in[5] ui_in[4] 0.023797f
C264 uio_oe[6] uio_oe[7] 0.023797f
C265 uo_out[0] uo_out[2] 0.013858f
C266 ui_in[0] X_TIMER.q_sr 0.021046f
C267 uo_out[0] uio_out[5] 0.013858f
C268 uio_out[7] uio_out[6] 0.023797f
C269 X_TIMER.X_COMP_P_TOP.latch_left ua[0] 0.533218f
C270 X_TIMER.X_COMP_P_TOP.out_left X_TIMER.X_SR_LATCH.IN_S 0.016125f
C271 ua[3] VGND 0.101433f
C272 ua[4] VGND 0.101433f
C273 ua[5] VGND 0.101909f
C274 ua[6] VGND 0.102993f
C275 ua[7] VGND 0.111838f
C276 ena VGND 0.073297f
C277 clk VGND 0.0487f
C278 rst_n VGND 0.04861f
C279 ui_in[1] VGND 0.040051f
C280 ui_in[2] VGND 0.040155f
C281 ui_in[3] VGND 0.040155f
C282 ui_in[4] VGND 0.040155f
C283 ui_in[5] VGND 0.040155f
C284 ui_in[6] VGND 0.040155f
C285 ui_in[7] VGND 0.040155f
C286 uio_in[0] VGND 0.040155f
C287 uio_in[1] VGND 0.040155f
C288 uio_in[2] VGND 0.040155f
C289 uio_in[3] VGND 0.040155f
C290 uio_in[4] VGND 0.040155f
C291 uio_in[5] VGND 0.040155f
C292 uio_in[6] VGND 0.040155f
C293 uio_in[7] VGND 0.040155f
C294 uo_out[1] VGND 0.03939f
C295 uo_out[2] VGND 0.03939f
C296 uo_out[3] VGND 0.03939f
C297 uo_out[4] VGND 0.03939f
C298 uo_out[5] VGND 0.03939f
C299 uo_out[6] VGND 0.03939f
C300 uo_out[7] VGND 0.03939f
C301 uio_out[0] VGND 0.03939f
C302 uio_out[1] VGND 0.03939f
C303 uio_out[2] VGND 0.03939f
C304 uio_out[3] VGND 0.03939f
C305 uio_out[4] VGND 0.03939f
C306 uio_out[5] VGND 0.03939f
C307 uio_out[6] VGND 0.03939f
C308 uio_out[7] VGND 0.03939f
C309 uio_oe[0] VGND 0.03939f
C310 uio_oe[1] VGND 0.03939f
C311 uio_oe[2] VGND 0.03939f
C312 uio_oe[3] VGND 0.03939f
C313 uio_oe[4] VGND 0.03939f
C314 uio_oe[5] VGND 0.03939f
C315 uio_oe[6] VGND 0.03939f
C316 uio_oe[7] VGND 0.073297f
C317 ua[2] VGND 21.234564f
C318 ua[1] VGND 29.932108f
C319 uo_out[0] VGND 26.68811f
C320 ui_in[0] VGND 41.601727f
C321 ua[0] VGND 31.993484f
C322 VPWR VGND 0.117201p
C323 X_TIMER.X_SR_LATCH.nand_0.drain_mna VGND 0.108562f
C324 X_TIMER.X_COMP_P_BOTTOM.latch_right VGND 7.51664f
C325 X_TIMER.X_COMP_P_BOTTOM.latch_left VGND 6.360844f
C326 X_TIMER.out_inv3 VGND 4.3233f
C327 a_1723_2994# VGND 0.023021f
C328 a_1347_2994# VGND 0.023021f
C329 X_TIMER.out_inv1 VGND 0.809774f
C330 X_TIMER.X_SR_LATCH.X_NOR_BOTTOM.IN_B VGND 0.488682f
C331 X_TIMER.qb_sr VGND 0.601493f
C332 X_TIMER.q_sr VGND 0.845576f
C333 X_TIMER.X_SR_LATCH.nand_0.IN_A VGND 0.587746f
C334 X_TIMER.X_COMP_P_BOTTOM.tail VGND 3.33693f
C335 X_TIMER.X_SR_LATCH.IN_S VGND 11.865175f
C336 X_TIMER.X_COMP_P_BOTTOM.out_left VGND 4.02347f
C337 X_TIMER.v0p6 VGND 2.29578f
C338 X_TIMER.v1p2 VGND 3.36574f
C339 X_TIMER.X_COMP_P_TOP.tail VGND 3.32219f
C340 X_TIMER.bias_p VGND 2.55084f
C341 X_TIMER.bias_1 VGND 1.57698f
C342 X_TIMER.bias_2 VGND 1.43453f
C343 X_TIMER.bias_3 VGND 1.65425f
C344 X_TIMER.X_COMP_P_TOP.latch_right VGND 6.586444f
C345 X_TIMER.X_COMP_P_TOP.out_left VGND 4.0365f
C346 X_TIMER.X_COMP_P_TOP.latch_left VGND 6.313573f
C347 X_TIMER.bias_n VGND 2.76281f
C348 ua[2].t1 VGND 0.129177f
C349 ua[2].t3 VGND 0.028175f
C350 ua[2].t0 VGND 0.028175f
C351 ua[2].n0 VGND 0.091167f
C352 ua[2].n1 VGND 0.497242f
C353 ua[2].t2 VGND 0.028175f
C354 ua[2].t4 VGND 0.028175f
C355 ua[2].n2 VGND 0.091167f
C356 ua[2].n3 VGND 0.393423f
C357 ua[2].n4 VGND 1.67706f
C358 X_TIMER.X_COMP_P_TOP.latch_left.t5 VGND 0.195314f
C359 X_TIMER.X_COMP_P_TOP.latch_left.t4 VGND 0.653259f
C360 X_TIMER.X_COMP_P_TOP.latch_left.t7 VGND 0.818972f
C361 X_TIMER.X_COMP_P_TOP.latch_left.t8 VGND 0.760557f
C362 X_TIMER.X_COMP_P_TOP.latch_left.n0 VGND 1.44598f
C363 X_TIMER.X_COMP_P_TOP.latch_left.n1 VGND 0.92801f
C364 X_TIMER.X_COMP_P_TOP.latch_left.n2 VGND 0.513842f
C365 X_TIMER.X_COMP_P_TOP.latch_left.t6 VGND 0.373955f
C366 X_TIMER.X_COMP_P_TOP.latch_left.t0 VGND 0.626969f
C367 X_TIMER.X_COMP_P_TOP.latch_left.t2 VGND 0.615096f
C368 X_TIMER.X_COMP_P_TOP.latch_left.n3 VGND 1.67064f
C369 X_TIMER.X_COMP_P_TOP.latch_left.n4 VGND 1.48416f
C370 X_TIMER.X_COMP_P_TOP.latch_left.n5 VGND 0.724094f
C371 X_TIMER.X_COMP_P_TOP.latch_left.t3 VGND 0.651869f
C372 X_TIMER.X_COMP_P_TOP.latch_left.t1 VGND 0.638869f
C373 X_TIMER.X_COMP_P_TOP.latch_left.n6 VGND 1.90364f
C374 X_TIMER.X_COMP_P_BOTTOM.out_left.n0 VGND 1.36437f
C375 X_TIMER.X_COMP_P_BOTTOM.out_left.n1 VGND 1.73513f
C376 X_TIMER.X_COMP_P_BOTTOM.out_left.t2 VGND 0.263818f
C377 X_TIMER.X_COMP_P_BOTTOM.out_left.t1 VGND 0.305396f
C378 X_TIMER.X_COMP_P_BOTTOM.out_left.t3 VGND 0.818674f
C379 X_TIMER.X_COMP_P_BOTTOM.out_left.t0 VGND 0.808807f
C380 X_TIMER.X_COMP_P_BOTTOM.latch_left.t3 VGND 0.651869f
C381 X_TIMER.X_COMP_P_BOTTOM.latch_left.t4 VGND 0.638869f
C382 X_TIMER.X_COMP_P_BOTTOM.latch_left.n0 VGND 1.90364f
C383 X_TIMER.X_COMP_P_BOTTOM.latch_left.t2 VGND 0.195313f
C384 X_TIMER.X_COMP_P_BOTTOM.latch_left.t1 VGND 0.653259f
C385 X_TIMER.X_COMP_P_BOTTOM.latch_left.t7 VGND 0.818972f
C386 X_TIMER.X_COMP_P_BOTTOM.latch_left.t8 VGND 0.760557f
C387 X_TIMER.X_COMP_P_BOTTOM.latch_left.n1 VGND 1.44598f
C388 X_TIMER.X_COMP_P_BOTTOM.latch_left.n2 VGND 0.92801f
C389 X_TIMER.X_COMP_P_BOTTOM.latch_left.n3 VGND 0.513842f
C390 X_TIMER.X_COMP_P_BOTTOM.latch_left.t5 VGND 0.626969f
C391 X_TIMER.X_COMP_P_BOTTOM.latch_left.t6 VGND 0.615096f
C392 X_TIMER.X_COMP_P_BOTTOM.latch_left.n4 VGND 1.67064f
C393 X_TIMER.X_COMP_P_BOTTOM.latch_left.t0 VGND 0.373955f
C394 X_TIMER.X_COMP_P_BOTTOM.latch_left.n5 VGND 1.48416f
C395 X_TIMER.X_COMP_P_BOTTOM.latch_left.n6 VGND 0.724094f
C396 ua[1].t3 VGND 0.716239f
C397 ua[1].t2 VGND 0.715763f
C398 ua[1].n0 VGND 0.63389f
C399 ua[1].n1 VGND 0.941039f
C400 ua[1].t1 VGND 0.531641f
C401 ua[1].t0 VGND 0.530955f
C402 ua[1].n2 VGND 0.773909f
C403 ua[1].n3 VGND 0.867187f
C404 ua[1].n4 VGND 0.455563f
C405 ui_in[0].t0 VGND 0.045708f
C406 ui_in[0].t1 VGND 0.02013f
C407 ui_in[0].n0 VGND 0.048111f
C408 ui_in[0].n1 VGND 0.007175f
C409 ui_in[0].n2 VGND 0.072481f
C410 X_TIMER.X_SR_LATCH.inv_0.vin VGND 2.01547f
C411 X_TIMER.X_SR_LATCH.IN_R.t3 VGND 0.034688f
C412 X_TIMER.X_SR_LATCH.IN_R.t2 VGND 0.034173f
C413 X_TIMER.X_SR_LATCH.IN_R.t1 VGND 0.41453f
C414 X_TIMER.X_SR_LATCH.IN_R.n0 VGND 3.09821f
C415 X_TIMER.X_SR_LATCH.IN_R.t0 VGND 0.533219f
C416 X_TIMER.X_COMP_P_TOP.vout VGND 1.66972f
C417 X_TIMER.X_COMP_P_TOP.out_left.n0 VGND 1.36437f
C418 X_TIMER.X_COMP_P_TOP.out_left.n1 VGND 1.73513f
C419 X_TIMER.X_COMP_P_TOP.out_left.t2 VGND 0.263818f
C420 X_TIMER.X_COMP_P_TOP.out_left.t1 VGND 0.305396f
C421 X_TIMER.X_COMP_P_TOP.out_left.t3 VGND 0.818674f
C422 X_TIMER.X_COMP_P_TOP.out_left.t0 VGND 0.808807f
C423 X_TIMER.X_SR_LATCH.IN_S.t3 VGND 0.028431f
C424 X_TIMER.X_SR_LATCH.IN_S.t2 VGND 0.012521f
C425 X_TIMER.X_SR_LATCH.IN_S.n0 VGND 0.029852f
C426 X_TIMER.X_SR_LATCH.IN_S.n1 VGND 0.635801f
C427 X_TIMER.X_SR_LATCH.IN_S.t1 VGND 0.140783f
C428 X_TIMER.X_SR_LATCH.IN_S.n2 VGND 1.20414f
C429 X_TIMER.X_SR_LATCH.IN_S.t0 VGND 0.299496f
C430 X_TIMER.X_COMP_P_BOTTOM.tail.t6 VGND 1.24327f
C431 X_TIMER.X_COMP_P_BOTTOM.tail.t3 VGND 1.23117f
C432 X_TIMER.X_COMP_P_BOTTOM.tail.n0 VGND 3.22105f
C433 X_TIMER.X_COMP_P_BOTTOM.tail.t7 VGND 1.2318f
C434 X_TIMER.X_COMP_P_BOTTOM.tail.n1 VGND 1.67554f
C435 X_TIMER.X_COMP_P_BOTTOM.tail.t1 VGND 1.23124f
C436 X_TIMER.X_COMP_P_BOTTOM.tail.n2 VGND 1.66379f
C437 X_TIMER.X_COMP_P_BOTTOM.tail.t8 VGND 0.996939f
C438 X_TIMER.X_COMP_P_BOTTOM.tail.t2 VGND 1.24361f
C439 X_TIMER.X_COMP_P_BOTTOM.tail.t4 VGND 1.23219f
C440 X_TIMER.X_COMP_P_BOTTOM.tail.n3 VGND 3.21408f
C441 X_TIMER.X_COMP_P_BOTTOM.tail.t0 VGND 1.23219f
C442 X_TIMER.X_COMP_P_BOTTOM.tail.n4 VGND 1.67418f
C443 X_TIMER.X_COMP_P_BOTTOM.tail.t5 VGND 1.23219f
C444 X_TIMER.X_COMP_P_BOTTOM.tail.n5 VGND 1.69154f
C445 X_TIMER.X_COMP_P_TOP.latch_right.n0 VGND 0.641993f
C446 X_TIMER.X_COMP_P_TOP.latch_right.n1 VGND 1.16334f
C447 X_TIMER.X_COMP_P_TOP.latch_right.t2 VGND 0.248107f
C448 X_TIMER.X_COMP_P_TOP.latch_right.t7 VGND 1.04034f
C449 X_TIMER.X_COMP_P_TOP.latch_right.t8 VGND 0.966138f
C450 X_TIMER.X_COMP_P_TOP.latch_right.n2 VGND 1.82161f
C451 X_TIMER.X_COMP_P_TOP.latch_right.t1 VGND 0.82985f
C452 X_TIMER.X_COMP_P_TOP.latch_right.t3 VGND 0.80961f
C453 X_TIMER.X_COMP_P_TOP.latch_right.t6 VGND 0.795083f
C454 X_TIMER.X_COMP_P_TOP.latch_right.n3 VGND 2.26592f
C455 X_TIMER.X_COMP_P_TOP.latch_right.t0 VGND 0.46252f
C456 X_TIMER.X_COMP_P_TOP.latch_right.t5 VGND 0.79635f
C457 X_TIMER.X_COMP_P_TOP.latch_right.t4 VGND 0.781068f
C458 X_TIMER.X_COMP_P_TOP.latch_right.n4 VGND 2.10739f
C459 X_TIMER.X_COMP_P_TOP.latch_right.n5 VGND 1.90069f
C460 X_TIMER.X_COMP_P_TOP.latch_right.n6 VGND 0.90098f
C461 X_TIMER.X_COMP_P_TOP.tail.n0 VGND 3.17699f
C462 X_TIMER.X_COMP_P_TOP.tail.n1 VGND 3.32689f
C463 X_TIMER.X_COMP_P_TOP.tail.n2 VGND 3.18388f
C464 X_TIMER.X_COMP_P_TOP.tail.n3 VGND 3.30081f
C465 X_TIMER.X_COMP_P_TOP.tail.t0 VGND 1.22892f
C466 X_TIMER.X_COMP_P_TOP.tail.t8 VGND 1.21696f
C467 X_TIMER.X_COMP_P_TOP.tail.t2 VGND 1.21758f
C468 X_TIMER.X_COMP_P_TOP.tail.t7 VGND 1.21703f
C469 X_TIMER.X_COMP_P_TOP.tail.t4 VGND 0.985436f
C470 X_TIMER.X_COMP_P_TOP.tail.t5 VGND 1.22926f
C471 X_TIMER.X_COMP_P_TOP.tail.t3 VGND 1.21797f
C472 X_TIMER.X_COMP_P_TOP.tail.t6 VGND 1.21797f
C473 X_TIMER.X_COMP_P_TOP.tail.t1 VGND 1.21797f
C474 ua[0].t0 VGND 0.561754f
C475 ua[0].t3 VGND 0.561381f
C476 ua[0].n0 VGND 0.75427f
C477 ua[0].n1 VGND 0.590521f
C478 ua[0].t2 VGND 0.417497f
C479 ua[0].n2 VGND 0.679183f
C480 ua[0].t1 VGND 0.416963f
C481 ua[0].n3 VGND 0.667757f
C482 ua[0].n4 VGND 0.316491f
C483 X_TIMER.X_COMP_P_BOTTOM.latch_right.n0 VGND 4.0306f
C484 X_TIMER.X_COMP_P_BOTTOM.latch_right.n1 VGND 0.645599f
C485 X_TIMER.X_COMP_P_BOTTOM.latch_right.n2 VGND 1.16988f
C486 X_TIMER.X_COMP_P_BOTTOM.latch_right.t1 VGND 0.814158f
C487 X_TIMER.X_COMP_P_BOTTOM.latch_right.t3 VGND 0.79955f
C488 X_TIMER.X_COMP_P_BOTTOM.latch_right.n3 VGND 2.27865f
C489 X_TIMER.X_COMP_P_BOTTOM.latch_right.t0 VGND 0.800824f
C490 X_TIMER.X_COMP_P_BOTTOM.latch_right.t2 VGND 0.785456f
C491 X_TIMER.X_COMP_P_BOTTOM.latch_right.t4 VGND 0.465119f
C492 X_TIMER.X_COMP_P_BOTTOM.latch_right.t6 VGND 0.249501f
C493 X_TIMER.X_COMP_P_BOTTOM.latch_right.t7 VGND 1.04619f
C494 X_TIMER.X_COMP_P_BOTTOM.latch_right.t8 VGND 0.971566f
C495 X_TIMER.X_COMP_P_BOTTOM.latch_right.n4 VGND 1.83184f
C496 X_TIMER.X_COMP_P_BOTTOM.latch_right.t5 VGND 0.834512f
C497 VPWR.n0 VGND 1.41928f
C498 VPWR.n1 VGND 0.218773f
C499 VPWR.n2 VGND 0.291021f
C500 VPWR.n3 VGND 0.123558f
C501 VPWR.t36 VGND 0.100664f
C502 VPWR.n4 VGND 0.115224f
C503 VPWR.n5 VGND 0.04621f
C504 VPWR.n6 VGND 0.04621f
C505 VPWR.t37 VGND 2.36013f
C506 VPWR.n7 VGND 0.055003f
C507 VPWR.n8 VGND 0.118525f
C508 VPWR.n9 VGND 0.128123f
C509 VPWR.n10 VGND 0.045202f
C510 VPWR.n11 VGND 0.045202f
C511 VPWR.n12 VGND 0.045202f
C512 VPWR.t39 VGND 2.41513f
C513 VPWR.n13 VGND 0.058208f
C514 VPWR.n14 VGND 0.035101f
C515 VPWR.n15 VGND 0.032504f
C516 VPWR.n16 VGND 0.032456f
C517 VPWR.n17 VGND 0.010511f
C518 VPWR.n18 VGND 0.230437f
C519 VPWR.n19 VGND 0.521382f
C520 VPWR.n20 VGND 1.76455f
C521 VPWR.n21 VGND 0.488757f
C522 VPWR.n22 VGND 0.123558f
C523 VPWR.n23 VGND 0.045463f
C524 VPWR.n24 VGND 0.007352f
C525 VPWR.n25 VGND 0.128123f
C526 VPWR.n26 VGND 0.035101f
C527 VPWR.n27 VGND 0.063764f
C528 VPWR.n28 VGND 0.233178f
C529 VPWR.n29 VGND 1.97011f
C530 VPWR.n30 VGND 2.27195f
C531 VPWR.n31 VGND 0.117941f
C532 VPWR.n32 VGND 0.035211f
C533 VPWR.n33 VGND 0.41082f
C534 VPWR.n34 VGND 0.041691f
C535 VPWR.n35 VGND 0.006425f
C536 VPWR.n36 VGND 0.045373f
C537 VPWR.n37 VGND 0.417523f
C538 VPWR.n38 VGND 0.045463f
C539 VPWR.n39 VGND 0.006425f
C540 VPWR.n40 VGND 0.041691f
C541 VPWR.n41 VGND 0.045373f
C542 VPWR.n42 VGND 0.016493f
C543 VPWR.n43 VGND 0.072309f
C544 VPWR.n44 VGND 0.118525f
C545 VPWR.n45 VGND 0.122507f
C546 VPWR.n46 VGND 0.010001f
C547 VPWR.n47 VGND 0.045202f
C548 VPWR.n48 VGND 0.021297f
C549 VPWR.n49 VGND 0.398219f
C550 VPWR.t19 VGND 0.417523f
C551 VPWR.n50 VGND 0.054532f
C552 VPWR.n51 VGND 0.054532f
C553 VPWR.n52 VGND 0.032456f
C554 VPWR.n53 VGND 0.015713f
C555 VPWR.n54 VGND 0.019405f
C556 VPWR.n55 VGND 0.032504f
C557 VPWR.n56 VGND 0.06381f
C558 VPWR.n57 VGND 0.035201f
C559 VPWR.n58 VGND 2.27439f
C560 VPWR.n59 VGND 0.04621f
C561 VPWR.n60 VGND 1.8601f
C562 VPWR.t12 VGND 0.010001f
C563 VPWR.t1 VGND 0.422523f
C564 VPWR.t21 VGND 0.422523f
C565 VPWR.n61 VGND 0.054532f
C566 VPWR.n62 VGND 0.007352f
C567 VPWR.n63 VGND 0.058208f
C568 VPWR.n64 VGND 0.054532f
C569 VPWR.t25 VGND 2.36013f
C570 VPWR.n65 VGND 0.035206f
C571 VPWR.n66 VGND 0.041701f
C572 VPWR.n67 VGND 0.045357f
C573 VPWR.n68 VGND 0.045357f
C574 VPWR.n69 VGND 0.054083f
C575 VPWR.n70 VGND 0.242944f
C576 VPWR.n71 VGND 0.021297f
C577 VPWR.n72 VGND 0.398219f
C578 VPWR.n73 VGND 0.72941f
C579 VPWR.n74 VGND 0.2312f
C580 VPWR.n75 VGND 0.023513f
C581 VPWR.n76 VGND 1.8601f
C582 VPWR.n77 VGND 0.847547f
C583 VPWR.n78 VGND 0.023539f
C584 VPWR.n79 VGND 0.2312f
C585 VPWR.n80 VGND 0.72941f
C586 VPWR.n81 VGND 0.242944f
C587 VPWR.n82 VGND 0.117699f
C588 VPWR.n83 VGND 0.126979f
C589 VPWR.n84 VGND 0.016493f
C590 VPWR.n85 VGND 0.045202f
C591 VPWR.n86 VGND 0.041701f
C592 VPWR.n87 VGND 0.045357f
C593 VPWR.n88 VGND 0.122507f
C594 VPWR.n89 VGND 0.045357f
C595 VPWR.n90 VGND 0.045202f
C596 VPWR.n91 VGND 0.045373f
C597 VPWR.n92 VGND 0.054312f
C598 VPWR.n93 VGND 0.244292f
C599 VPWR.n94 VGND 0.746792f
C600 VPWR.n95 VGND 0.41082f
C601 VPWR.n96 VGND 0.04621f
C602 VPWR.n97 VGND 0.017501f
C603 VPWR.t0 VGND 0.017501f
C604 VPWR.t11 VGND 0.010001f
C605 VPWR.n98 VGND 0.010001f
C606 VPWR.n99 VGND 0.045373f
C607 VPWR.n100 VGND 0.072476f
C608 VPWR.n101 VGND 0.244292f
C609 VPWR.n102 VGND 0.746792f
C610 VPWR.n103 VGND 0.233178f
C611 VPWR.n104 VGND 0.023523f
C612 VPWR.n105 VGND 0.850047f
C613 VPWR.n106 VGND 1.97011f
C614 VPWR.n107 VGND 0.023513f
C615 VPWR.n108 VGND 0.035206f
C616 VPWR.n109 VGND 0.117941f
C617 VPWR.n110 VGND 0.115224f
C618 VPWR.t38 VGND 0.100664f
C619 VPWR.n111 VGND 0.11939f
C620 VPWR.n112 VGND 0.057439f
C621 VPWR.n113 VGND 0.219476f
C622 VPWR.n114 VGND 0.04621f
C623 VPWR.n115 VGND 0.045463f
C624 VPWR.n116 VGND 0.045463f
C625 VPWR.n117 VGND 0.045463f
C626 VPWR.n118 VGND 0.399474f
C627 VPWR.t33 VGND 0.674428f
C628 VPWR.n121 VGND 0.399474f
C629 VPWR.n122 VGND 0.04621f
C630 VPWR.n123 VGND 0.045463f
C631 VPWR.t34 VGND 0.101779f
C632 VPWR.n124 VGND 0.465931f
C633 VPWR.n125 VGND 1.48785f
C634 VPWR.n126 VGND 1.12665f
C635 VPWR.n127 VGND 0.334992f
C636 VPWR.n128 VGND 0.238515f
C637 VPWR.t26 VGND 0.081463f
C638 VPWR.n129 VGND 0.146815f
C639 VPWR.t22 VGND 0.081463f
C640 VPWR.n130 VGND 0.194599f
C641 VPWR.n131 VGND 0.633984f
C642 VPWR.n132 VGND 0.275661f
C643 VPWR.n133 VGND 2.3656f
C644 VPWR.n134 VGND 0.410119f
C645 VPWR.n135 VGND 0.289936f
C646 VPWR.n136 VGND 0.099531f
C647 VPWR.n137 VGND 0.266767f
C648 VPWR.t20 VGND 0.081463f
C649 VPWR.n138 VGND 0.194599f
C650 VPWR.t40 VGND 0.081463f
C651 VPWR.n139 VGND 0.194599f
C652 VPWR.n140 VGND 0.40846f
C653 VPWR.n141 VGND 0.156625f
C654 VPWR.n142 VGND 0.011008f
C655 VPWR.n143 VGND 0.015713f
C656 VPWR.n144 VGND 0.019405f
C657 VPWR.n145 VGND 0.007352f
C658 VPWR.n146 VGND 0.007352f
C659 VPWR.n147 VGND 2.41513f
C660 VPWR.n148 VGND 0.016493f
C661 VPWR.n149 VGND 0.016493f
C662 VPWR.n150 VGND 0.126979f
C663 VPWR.n151 VGND 0.117699f
C664 VPWR.n152 VGND 0.045463f
C665 VPWR.t35 VGND 0.055003f
C666 VPWR.n153 VGND 0.045463f
C667 VPWR.n154 VGND 0.11939f
C668 VPWR.n155 VGND 0.057698f
C669 VPWR.n156 VGND 0.488847f
C670 VPWR.n157 VGND 1.1651f
C671 VPWR.t30 VGND 0.010225f
C672 VPWR.n158 VGND 0.020197f
C673 VPWR.n159 VGND 0.008556f
C674 VPWR.n160 VGND 0.00854f
C675 VPWR.n161 VGND 0.006269f
C676 VPWR.n162 VGND 0.012344f
C677 VPWR.t8 VGND 0.163045f
C678 VPWR.n163 VGND 0.008556f
C679 VPWR.n164 VGND 0.008556f
C680 VPWR.t5 VGND 0.010225f
C681 VPWR.t7 VGND 0.010225f
C682 VPWR.t3 VGND 0.010225f
C683 VPWR.n165 VGND 0.026603f
C684 VPWR.n166 VGND 0.008995f
C685 VPWR.n167 VGND 0.007661f
C686 VPWR.t2 VGND 0.170778f
C687 VPWR.t4 VGND 0.164823f
C688 VPWR.t6 VGND 0.164823f
C689 VPWR.n168 VGND 0.008556f
C690 VPWR.n169 VGND 0.008556f
C691 VPWR.n170 VGND 0.006295f
C692 VPWR.n171 VGND 0.020197f
C693 VPWR.n172 VGND 0.006295f
C694 VPWR.n173 VGND 0.020197f
C695 VPWR.t9 VGND 0.010225f
C696 VPWR.t32 VGND 0.010225f
C697 VPWR.n174 VGND 0.020197f
C698 VPWR.n175 VGND 0.006295f
C699 VPWR.n176 VGND 0.020197f
C700 VPWR.n177 VGND 0.006295f
C701 VPWR.n178 VGND 0.008556f
C702 VPWR.n179 VGND 0.008556f
C703 VPWR.n180 VGND 0.008556f
C704 VPWR.t31 VGND 0.164823f
C705 VPWR.t29 VGND 0.164511f
C706 VPWR.t15 VGND 0.102797f
C707 VPWR.n181 VGND 0.011251f
C708 VPWR.t44 VGND 0.020536f
C709 VPWR.t18 VGND 0.010225f
C710 VPWR.n182 VGND 0.020197f
C711 VPWR.n183 VGND 0.017565f
C712 VPWR.n184 VGND 0.038127f
C713 VPWR.t16 VGND 0.020536f
C714 VPWR.t14 VGND 0.010225f
C715 VPWR.n185 VGND 0.019743f
C716 VPWR.t23 VGND 0.101112f
C717 VPWR.n186 VGND 0.027575f
C718 VPWR.t41 VGND 0.1009f
C719 VPWR.t13 VGND 0.174225f
C720 VPWR.n187 VGND 0.00906f
C721 VPWR.n188 VGND 0.01417f
C722 VPWR.t24 VGND 0.005549f
C723 VPWR.t42 VGND 0.005549f
C724 VPWR.n189 VGND 0.016924f
C725 VPWR.n190 VGND 0.018639f
C726 VPWR.n191 VGND 0.008065f
C727 VPWR.n192 VGND 0.038127f
C728 VPWR.n193 VGND 0.017748f
C729 VPWR.n194 VGND 0.013012f
C730 VPWR.n195 VGND 0.027574f
C731 VPWR.t27 VGND 0.103093f
C732 VPWR.t43 VGND 0.104973f
C733 VPWR.n196 VGND 0.027574f
C734 VPWR.t10 VGND 0.103093f
C735 VPWR.t17 VGND 0.172345f
C736 VPWR.n197 VGND 0.009604f
C737 VPWR.n198 VGND 0.008849f
C738 VPWR.n199 VGND 0.00854f
C739 VPWR.n200 VGND 0.005583f
C740 VPWR.n201 VGND 0.094227f
C741 VPWR.n202 VGND 1.36629f
C742 VPWR.n203 VGND 12.834599f
C743 uo_out[0].t5 VGND 0.041612f
C744 uo_out[0].t9 VGND 0.041612f
C745 uo_out[0].t10 VGND 0.041612f
C746 uo_out[0].t6 VGND 0.041612f
C747 uo_out[0].t1 VGND 0.061878f
C748 uo_out[0].t3 VGND 0.060757f
C749 uo_out[0].t2 VGND 0.061878f
C750 uo_out[0].t0 VGND 0.060757f
C751 uo_out[0].n0 VGND 0.363072f
C752 uo_out[0].n1 VGND 0.383058f
C753 uo_out[0].t4 VGND 0.040335f
C754 uo_out[0].n2 VGND 0.082139f
C755 uo_out[0].n3 VGND 0.171418f
C756 uo_out[0].t8 VGND 0.040994f
C757 uo_out[0].n4 VGND 0.229344f
C758 uo_out[0].t7 VGND 0.040994f
C759 uo_out[0].n5 VGND 0.229344f
C760 uo_out[0].t11 VGND 0.040994f
C761 uo_out[0].n6 VGND 1.66329f
C762 uo_out[0].n7 VGND 9.82069f
.ends

