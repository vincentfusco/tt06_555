magic
tech sky130A
magscale 1 2
timestamp 1710860643
<< error_p >>
rect -77 1181 -19 1187
rect -77 1147 -65 1181
rect -77 1141 -19 1147
rect 19 71 77 77
rect 19 37 31 71
rect 19 31 77 37
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 19 -77 77 -71
rect -77 -1147 -19 -1141
rect -77 -1181 -65 -1147
rect -77 -1187 -19 -1181
<< pwell >>
rect -263 -1319 263 1319
<< nmos >>
rect -63 109 -33 1109
rect 33 109 63 1109
rect -63 -1109 -33 -109
rect 33 -1109 63 -109
<< ndiff >>
rect -125 1097 -63 1109
rect -125 121 -113 1097
rect -79 121 -63 1097
rect -125 109 -63 121
rect -33 1097 33 1109
rect -33 121 -17 1097
rect 17 121 33 1097
rect -33 109 33 121
rect 63 1097 125 1109
rect 63 121 79 1097
rect 113 121 125 1097
rect 63 109 125 121
rect -125 -121 -63 -109
rect -125 -1097 -113 -121
rect -79 -1097 -63 -121
rect -125 -1109 -63 -1097
rect -33 -121 33 -109
rect -33 -1097 -17 -121
rect 17 -1097 33 -121
rect -33 -1109 33 -1097
rect 63 -121 125 -109
rect 63 -1097 79 -121
rect 113 -1097 125 -121
rect 63 -1109 125 -1097
<< ndiffc >>
rect -113 121 -79 1097
rect -17 121 17 1097
rect 79 121 113 1097
rect -113 -1097 -79 -121
rect -17 -1097 17 -121
rect 79 -1097 113 -121
<< psubdiff >>
rect -227 1249 -131 1283
rect 131 1249 227 1283
rect -227 1187 -193 1249
rect 193 1187 227 1249
rect -227 -1249 -193 -1187
rect 193 -1249 227 -1187
rect -227 -1283 -131 -1249
rect 131 -1283 227 -1249
<< psubdiffcont >>
rect -131 1249 131 1283
rect -227 -1187 -193 1187
rect 193 -1187 227 1187
rect -131 -1283 131 -1249
<< poly >>
rect -81 1181 -15 1197
rect -81 1147 -65 1181
rect -31 1147 -15 1181
rect -81 1131 -15 1147
rect -63 1109 -33 1131
rect 33 1109 63 1135
rect -63 83 -33 109
rect 33 87 63 109
rect 15 71 81 87
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 33 -109 63 -87
rect -63 -1131 -33 -1109
rect -81 -1147 -15 -1131
rect 33 -1135 63 -1109
rect -81 -1181 -65 -1147
rect -31 -1181 -15 -1147
rect -81 -1197 -15 -1181
<< polycont >>
rect -65 1147 -31 1181
rect 31 37 65 71
rect 31 -71 65 -37
rect -65 -1181 -31 -1147
<< locali >>
rect -227 1249 -131 1283
rect 131 1249 227 1283
rect -227 1187 -193 1249
rect 193 1187 227 1249
rect -81 1147 -65 1181
rect -31 1147 -15 1181
rect -113 1097 -79 1113
rect -113 105 -79 121
rect -17 1097 17 1113
rect -17 105 17 121
rect 79 1097 113 1113
rect 79 105 113 121
rect 15 37 31 71
rect 65 37 81 71
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -113 -121 -79 -105
rect -113 -1113 -79 -1097
rect -17 -121 17 -105
rect -17 -1113 17 -1097
rect 79 -121 113 -105
rect 79 -1113 113 -1097
rect -81 -1181 -65 -1147
rect -31 -1181 -15 -1147
rect -227 -1249 -193 -1187
rect 193 -1249 227 -1187
rect -227 -1283 -131 -1249
rect 131 -1283 227 -1249
<< viali >>
rect -65 1147 -31 1181
rect -113 121 -79 1097
rect -17 121 17 1097
rect 79 121 113 1097
rect 31 37 65 71
rect 31 -71 65 -37
rect -113 -1097 -79 -121
rect -17 -1097 17 -121
rect 79 -1097 113 -121
rect -65 -1181 -31 -1147
<< metal1 >>
rect -77 1181 -19 1187
rect -77 1147 -65 1181
rect -31 1147 -19 1181
rect -77 1141 -19 1147
rect -119 1097 -73 1109
rect -119 121 -113 1097
rect -79 121 -73 1097
rect -119 109 -73 121
rect -23 1097 23 1109
rect -23 121 -17 1097
rect 17 121 23 1097
rect -23 109 23 121
rect 73 1097 119 1109
rect 73 121 79 1097
rect 113 121 119 1097
rect 73 109 119 121
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect -119 -121 -73 -109
rect -119 -1097 -113 -121
rect -79 -1097 -73 -121
rect -119 -1109 -73 -1097
rect -23 -121 23 -109
rect -23 -1097 -17 -121
rect 17 -1097 23 -121
rect -23 -1109 23 -1097
rect 73 -121 119 -109
rect 73 -1097 79 -121
rect 113 -1097 119 -121
rect 73 -1109 119 -1097
rect -77 -1147 -19 -1141
rect -77 -1181 -65 -1147
rect -31 -1181 -19 -1147
rect -77 -1187 -19 -1181
<< properties >>
string FIXED_BBOX -210 -1266 210 1266
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
