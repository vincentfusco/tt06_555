magic
tech sky130A
magscale 1 2
timestamp 1711053111
<< checkpaint >>
rect 3278 3219 6390 3272
rect 3278 -1286 6929 3219
rect 3817 -1339 6929 -1286
<< error_s >>
rect 338 9623 373 9657
rect 339 9604 373 9623
rect 147 9555 209 9561
rect 147 9521 159 9555
rect 147 9515 209 9521
rect 147 7427 209 7433
rect 147 7393 159 7427
rect 147 7387 209 7393
rect 147 7319 209 7325
rect 147 7285 159 7319
rect 147 7279 209 7285
rect 147 5191 209 5197
rect 147 5157 159 5191
rect 147 5151 209 5157
rect 147 5083 209 5089
rect 147 5049 159 5083
rect 147 5043 209 5049
rect 147 2955 209 2961
rect 147 2921 159 2955
rect 147 2915 209 2921
rect 147 2847 209 2853
rect 147 2813 159 2847
rect 147 2807 209 2813
rect 147 719 209 725
rect 147 685 159 719
rect 147 679 209 685
rect 358 583 373 9604
rect 392 9570 427 9604
rect 392 583 426 9570
rect 556 9502 618 9508
rect 556 9468 568 9502
rect 556 9462 618 9468
rect 556 7374 618 7380
rect 556 7340 568 7374
rect 556 7334 618 7340
rect 556 7266 618 7272
rect 556 7232 568 7266
rect 556 7226 618 7232
rect 556 5138 618 5144
rect 556 5104 568 5138
rect 556 5098 618 5104
rect 556 5030 618 5036
rect 556 4996 568 5030
rect 556 4990 618 4996
rect 556 2902 618 2908
rect 556 2868 568 2902
rect 556 2862 618 2868
rect 556 2794 618 2800
rect 556 2760 568 2794
rect 556 2754 618 2760
rect 1374 1794 1826 1826
rect 1374 1760 1826 1772
rect 2957 1734 2991 1752
rect 748 1661 782 1679
rect 748 1625 818 1661
rect 765 1591 836 1625
rect 556 666 618 672
rect 556 632 568 666
rect 556 626 618 632
rect 392 549 407 583
rect 765 530 835 1591
rect 765 494 818 530
rect 1306 477 1321 1625
rect 1340 477 1374 1676
rect 2452 1664 2904 1696
rect 2452 1630 2904 1642
rect 1826 1495 1860 1549
rect 1340 443 1355 477
rect 1845 400 1860 1495
rect 1879 1461 1914 1495
rect 1879 400 1913 1461
rect 1879 366 1894 400
rect 2384 347 2399 1495
rect 2418 347 2452 1546
rect 2418 313 2433 347
rect 2921 270 2991 1734
rect 3443 1604 3477 1622
rect 3443 1568 3513 1604
rect 3460 1566 3531 1568
rect 3460 1545 3982 1566
rect 3460 1534 4016 1545
rect 3460 1512 3530 1534
rect 3982 1512 4016 1534
rect 4574 1527 4608 1545
rect 3460 1500 4016 1512
rect 3460 1478 3531 1500
rect 3981 1491 4016 1500
rect 2921 234 2974 270
rect 3460 217 3530 1478
rect 3460 181 3513 217
rect 4001 140 4016 1491
rect 4035 1489 4070 1491
rect 4035 1457 4521 1489
rect 4035 1435 4069 1457
rect 4035 1423 4521 1435
rect 4035 1401 4070 1423
rect 4035 140 4069 1401
rect 4035 106 4050 140
rect 4538 63 4608 1527
rect 4538 27 4591 63
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_cs_left
timestamp 1711041810
transform 1 0 1600 0 1 1098
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_cs_right1
timestamp 1711041810
transform 1 0 2678 0 1 968
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XMn_diode_left1
timestamp 1711036998
transform 1 0 1061 0 1 1051
box -296 -610 296 610
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XMn_diode_right
timestamp 1711036998
transform 1 0 2139 0 1 921
box -296 -610 296 610
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_out_left
timestamp 1711041810
transform 1 0 4295 0 1 761
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_out_right
timestamp 1711041810
transform 1 0 3756 0 1 838
box -296 -734 296 766
use sky130_fd_pr__pfet_01v8_lvt_5VNMZ8  XMp_diode_left1
timestamp 1711036998
transform 1 0 4834 0 1 993
box -296 -1019 296 1019
use sky130_fd_pr__pfet_01v8_lvt_ERPZ26  XMp_inn1
timestamp 1711036998
transform 1 0 178 0 1 5120
box -231 -4573 231 4573
use sky130_fd_pr__pfet_01v8_lvt_ERPZ26  XMp_inp1
timestamp 1711036998
transform 1 0 587 0 1 5067
box -231 -4573 231 4573
use sky130_fd_pr__pfet_01v8_lvt_5VNMZ8  XMp_out
timestamp 1711036998
transform 1 0 5373 0 1 940
box -296 -1019 296 1019
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_tail
timestamp 1711036998
transform 1 0 3217 0 1 1400
box -296 -1219 296 1219
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 vinp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 vinn
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vbias_p
port 5 nsew
<< end >>
