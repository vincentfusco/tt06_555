magic
tech sky130A
magscale 1 2
timestamp 1711736161
<< error_p >>
rect -31 10072 31 10078
rect -31 10038 -19 10072
rect -31 10032 31 10038
rect -31 -10038 31 -10032
rect -31 -10072 -19 -10038
rect -31 -10078 31 -10072
<< pwell >>
rect -231 -10210 231 10210
<< nmoslvt >>
rect -35 -10000 35 10000
<< ndiff >>
rect -93 9988 -35 10000
rect -93 -9988 -81 9988
rect -47 -9988 -35 9988
rect -93 -10000 -35 -9988
rect 35 9988 93 10000
rect 35 -9988 47 9988
rect 81 -9988 93 9988
rect 35 -10000 93 -9988
<< ndiffc >>
rect -81 -9988 -47 9988
rect 47 -9988 81 9988
<< psubdiff >>
rect -195 10140 -99 10174
rect 99 10140 195 10174
rect -195 10078 -161 10140
rect 161 10078 195 10140
rect -195 -10140 -161 -10078
rect 161 -10140 195 -10078
rect -195 -10174 -99 -10140
rect 99 -10174 195 -10140
<< psubdiffcont >>
rect -99 10140 99 10174
rect -195 -10078 -161 10078
rect 161 -10078 195 10078
rect -99 -10174 99 -10140
<< poly >>
rect -35 10072 35 10088
rect -35 10038 -19 10072
rect 19 10038 35 10072
rect -35 10000 35 10038
rect -35 -10038 35 -10000
rect -35 -10072 -19 -10038
rect 19 -10072 35 -10038
rect -35 -10088 35 -10072
<< polycont >>
rect -19 10038 19 10072
rect -19 -10072 19 -10038
<< locali >>
rect -195 10140 -99 10174
rect 99 10140 195 10174
rect -195 10078 -161 10140
rect 161 10078 195 10140
rect -35 10038 -19 10072
rect 19 10038 35 10072
rect -81 9988 -47 10004
rect -81 -10004 -47 -9988
rect 47 9988 81 10004
rect 47 -10004 81 -9988
rect -35 -10072 -19 -10038
rect 19 -10072 35 -10038
rect -195 -10140 -161 -10078
rect 161 -10140 195 -10078
rect -195 -10174 -99 -10140
rect 99 -10174 195 -10140
<< viali >>
rect -19 10038 19 10072
rect -81 -9988 -47 9988
rect 47 -9988 81 9988
rect -19 -10072 19 -10038
<< metal1 >>
rect -31 10072 31 10078
rect -31 10038 -19 10072
rect 19 10038 31 10072
rect -31 10032 31 10038
rect -87 9988 -41 10000
rect -87 -9988 -81 9988
rect -47 -9988 -41 9988
rect -87 -10000 -41 -9988
rect 41 9988 87 10000
rect 41 -9988 47 9988
rect 81 -9988 87 9988
rect 41 -10000 87 -9988
rect -31 -10038 31 -10032
rect -31 -10072 -19 -10038
rect 19 -10072 31 -10038
rect -31 -10078 31 -10072
<< properties >>
string FIXED_BBOX -178 -10157 178 10157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 100 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
