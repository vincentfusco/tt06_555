magic
tech sky130A
magscale 1 2
timestamp 1711036998
<< error_p >>
rect -31 4435 31 4441
rect -31 4401 -19 4435
rect -31 4395 31 4401
rect -31 2307 31 2313
rect -31 2273 -19 2307
rect -31 2267 31 2273
rect -31 2199 31 2205
rect -31 2165 -19 2199
rect -31 2159 31 2165
rect -31 71 31 77
rect -31 37 -19 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect -31 -77 31 -71
rect -31 -2165 31 -2159
rect -31 -2199 -19 -2165
rect -31 -2205 31 -2199
rect -31 -2273 31 -2267
rect -31 -2307 -19 -2273
rect -31 -2313 31 -2307
rect -31 -4401 31 -4395
rect -31 -4435 -19 -4401
rect -31 -4441 31 -4435
<< nwell >>
rect -231 -4573 231 4573
<< pmoslvt >>
rect -35 2354 35 4354
rect -35 118 35 2118
rect -35 -2118 35 -118
rect -35 -4354 35 -2354
<< pdiff >>
rect -93 4342 -35 4354
rect -93 2366 -81 4342
rect -47 2366 -35 4342
rect -93 2354 -35 2366
rect 35 4342 93 4354
rect 35 2366 47 4342
rect 81 2366 93 4342
rect 35 2354 93 2366
rect -93 2106 -35 2118
rect -93 130 -81 2106
rect -47 130 -35 2106
rect -93 118 -35 130
rect 35 2106 93 2118
rect 35 130 47 2106
rect 81 130 93 2106
rect 35 118 93 130
rect -93 -130 -35 -118
rect -93 -2106 -81 -130
rect -47 -2106 -35 -130
rect -93 -2118 -35 -2106
rect 35 -130 93 -118
rect 35 -2106 47 -130
rect 81 -2106 93 -130
rect 35 -2118 93 -2106
rect -93 -2366 -35 -2354
rect -93 -4342 -81 -2366
rect -47 -4342 -35 -2366
rect -93 -4354 -35 -4342
rect 35 -2366 93 -2354
rect 35 -4342 47 -2366
rect 81 -4342 93 -2366
rect 35 -4354 93 -4342
<< pdiffc >>
rect -81 2366 -47 4342
rect 47 2366 81 4342
rect -81 130 -47 2106
rect 47 130 81 2106
rect -81 -2106 -47 -130
rect 47 -2106 81 -130
rect -81 -4342 -47 -2366
rect 47 -4342 81 -2366
<< nsubdiff >>
rect -195 4503 -99 4537
rect 99 4503 195 4537
rect -195 4441 -161 4503
rect 161 4441 195 4503
rect -195 -4503 -161 -4441
rect 161 -4503 195 -4441
rect -195 -4537 -99 -4503
rect 99 -4537 195 -4503
<< nsubdiffcont >>
rect -99 4503 99 4537
rect -195 -4441 -161 4441
rect 161 -4441 195 4441
rect -99 -4537 99 -4503
<< poly >>
rect -35 4435 35 4451
rect -35 4401 -19 4435
rect 19 4401 35 4435
rect -35 4354 35 4401
rect -35 2307 35 2354
rect -35 2273 -19 2307
rect 19 2273 35 2307
rect -35 2257 35 2273
rect -35 2199 35 2215
rect -35 2165 -19 2199
rect 19 2165 35 2199
rect -35 2118 35 2165
rect -35 71 35 118
rect -35 37 -19 71
rect 19 37 35 71
rect -35 21 35 37
rect -35 -37 35 -21
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect -35 -118 35 -71
rect -35 -2165 35 -2118
rect -35 -2199 -19 -2165
rect 19 -2199 35 -2165
rect -35 -2215 35 -2199
rect -35 -2273 35 -2257
rect -35 -2307 -19 -2273
rect 19 -2307 35 -2273
rect -35 -2354 35 -2307
rect -35 -4401 35 -4354
rect -35 -4435 -19 -4401
rect 19 -4435 35 -4401
rect -35 -4451 35 -4435
<< polycont >>
rect -19 4401 19 4435
rect -19 2273 19 2307
rect -19 2165 19 2199
rect -19 37 19 71
rect -19 -71 19 -37
rect -19 -2199 19 -2165
rect -19 -2307 19 -2273
rect -19 -4435 19 -4401
<< locali >>
rect -195 4503 -99 4537
rect 99 4503 195 4537
rect -195 4441 -161 4503
rect 161 4441 195 4503
rect -35 4401 -19 4435
rect 19 4401 35 4435
rect -81 4342 -47 4358
rect -81 2350 -47 2366
rect 47 4342 81 4358
rect 47 2350 81 2366
rect -35 2273 -19 2307
rect 19 2273 35 2307
rect -35 2165 -19 2199
rect 19 2165 35 2199
rect -81 2106 -47 2122
rect -81 114 -47 130
rect 47 2106 81 2122
rect 47 114 81 130
rect -35 37 -19 71
rect 19 37 35 71
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect -81 -130 -47 -114
rect -81 -2122 -47 -2106
rect 47 -130 81 -114
rect 47 -2122 81 -2106
rect -35 -2199 -19 -2165
rect 19 -2199 35 -2165
rect -35 -2307 -19 -2273
rect 19 -2307 35 -2273
rect -81 -2366 -47 -2350
rect -81 -4358 -47 -4342
rect 47 -2366 81 -2350
rect 47 -4358 81 -4342
rect -35 -4435 -19 -4401
rect 19 -4435 35 -4401
rect -195 -4503 -161 -4441
rect 161 -4503 195 -4441
rect -195 -4537 -99 -4503
rect 99 -4537 195 -4503
<< viali >>
rect -19 4401 19 4435
rect -81 2366 -47 4342
rect 47 2366 81 4342
rect -19 2273 19 2307
rect -19 2165 19 2199
rect -81 130 -47 2106
rect 47 130 81 2106
rect -19 37 19 71
rect -19 -71 19 -37
rect -81 -2106 -47 -130
rect 47 -2106 81 -130
rect -19 -2199 19 -2165
rect -19 -2307 19 -2273
rect -81 -4342 -47 -2366
rect 47 -4342 81 -2366
rect -19 -4435 19 -4401
<< metal1 >>
rect -31 4435 31 4441
rect -31 4401 -19 4435
rect 19 4401 31 4435
rect -31 4395 31 4401
rect -87 4342 -41 4354
rect -87 2366 -81 4342
rect -47 2366 -41 4342
rect -87 2354 -41 2366
rect 41 4342 87 4354
rect 41 2366 47 4342
rect 81 2366 87 4342
rect 41 2354 87 2366
rect -31 2307 31 2313
rect -31 2273 -19 2307
rect 19 2273 31 2307
rect -31 2267 31 2273
rect -31 2199 31 2205
rect -31 2165 -19 2199
rect 19 2165 31 2199
rect -31 2159 31 2165
rect -87 2106 -41 2118
rect -87 130 -81 2106
rect -47 130 -41 2106
rect -87 118 -41 130
rect 41 2106 87 2118
rect 41 130 47 2106
rect 81 130 87 2106
rect 41 118 87 130
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect -87 -130 -41 -118
rect -87 -2106 -81 -130
rect -47 -2106 -41 -130
rect -87 -2118 -41 -2106
rect 41 -130 87 -118
rect 41 -2106 47 -130
rect 81 -2106 87 -130
rect 41 -2118 87 -2106
rect -31 -2165 31 -2159
rect -31 -2199 -19 -2165
rect 19 -2199 31 -2165
rect -31 -2205 31 -2199
rect -31 -2273 31 -2267
rect -31 -2307 -19 -2273
rect 19 -2307 31 -2273
rect -31 -2313 31 -2307
rect -87 -2366 -41 -2354
rect -87 -4342 -81 -2366
rect -47 -4342 -41 -2366
rect -87 -4354 -41 -4342
rect 41 -2366 87 -2354
rect 41 -4342 47 -2366
rect 81 -4342 87 -2366
rect 41 -4354 87 -4342
rect -31 -4401 31 -4395
rect -31 -4435 -19 -4401
rect 19 -4435 31 -4401
rect -31 -4441 31 -4435
<< properties >>
string FIXED_BBOX -178 -4520 178 4520
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 0.35 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
