magic
tech sky130A
magscale 1 2
timestamp 1711041017
<< error_p >>
rect -223 572 -161 578
rect -95 572 -33 578
rect 33 572 95 578
rect 161 572 223 578
rect -223 538 -211 572
rect -95 538 -83 572
rect 33 538 45 572
rect 161 538 173 572
rect -223 532 -161 538
rect -95 532 -33 538
rect 33 532 95 538
rect 161 532 223 538
rect -223 -538 -161 -532
rect -95 -538 -33 -532
rect 33 -538 95 -532
rect 161 -538 223 -532
rect -223 -572 -211 -538
rect -95 -572 -83 -538
rect 33 -572 45 -538
rect 161 -572 173 -538
rect -223 -578 -161 -572
rect -95 -578 -33 -572
rect 33 -578 95 -572
rect 161 -578 223 -572
<< pwell >>
rect -423 -710 423 710
<< nmoslvt >>
rect -227 -500 -157 500
rect -99 -500 -29 500
rect 29 -500 99 500
rect 157 -500 227 500
<< ndiff >>
rect -285 488 -227 500
rect -285 -488 -273 488
rect -239 -488 -227 488
rect -285 -500 -227 -488
rect -157 488 -99 500
rect -157 -488 -145 488
rect -111 -488 -99 488
rect -157 -500 -99 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 99 488 157 500
rect 99 -488 111 488
rect 145 -488 157 488
rect 99 -500 157 -488
rect 227 488 285 500
rect 227 -488 239 488
rect 273 -488 285 488
rect 227 -500 285 -488
<< ndiffc >>
rect -273 -488 -239 488
rect -145 -488 -111 488
rect -17 -488 17 488
rect 111 -488 145 488
rect 239 -488 273 488
<< psubdiff >>
rect -387 640 -291 674
rect 291 640 387 674
rect -387 -640 -353 640
rect 353 578 387 640
rect 353 -640 387 -578
rect -387 -674 -291 -640
rect 291 -674 387 -640
<< psubdiffcont >>
rect -291 640 291 674
rect 353 -578 387 578
rect -291 -674 291 -640
<< poly >>
rect -227 572 -157 588
rect -227 538 -211 572
rect -173 538 -157 572
rect -227 500 -157 538
rect -99 572 -29 588
rect -99 538 -83 572
rect -45 538 -29 572
rect -99 500 -29 538
rect 29 572 99 588
rect 29 538 45 572
rect 83 538 99 572
rect 29 500 99 538
rect 157 572 227 588
rect 157 538 173 572
rect 211 538 227 572
rect 157 500 227 538
rect -227 -538 -157 -500
rect -227 -572 -211 -538
rect -173 -572 -157 -538
rect -227 -588 -157 -572
rect -99 -538 -29 -500
rect -99 -572 -83 -538
rect -45 -572 -29 -538
rect -99 -588 -29 -572
rect 29 -538 99 -500
rect 29 -572 45 -538
rect 83 -572 99 -538
rect 29 -588 99 -572
rect 157 -538 227 -500
rect 157 -572 173 -538
rect 211 -572 227 -538
rect 157 -588 227 -572
<< polycont >>
rect -211 538 -173 572
rect -83 538 -45 572
rect 45 538 83 572
rect 173 538 211 572
rect -211 -572 -173 -538
rect -83 -572 -45 -538
rect 45 -572 83 -538
rect 173 -572 211 -538
<< locali >>
rect -387 640 -291 674
rect 291 640 387 674
rect -387 -640 -353 640
rect 353 578 387 640
rect -227 538 -211 572
rect -173 538 -157 572
rect -99 538 -83 572
rect -45 538 -29 572
rect 29 538 45 572
rect 83 538 99 572
rect 157 538 173 572
rect 211 538 227 572
rect -273 488 -239 504
rect -273 -504 -239 -488
rect -145 488 -111 504
rect -145 -504 -111 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 111 488 145 504
rect 111 -504 145 -488
rect 239 488 273 504
rect 239 -504 273 -488
rect -227 -572 -211 -538
rect -173 -572 -157 -538
rect -99 -572 -83 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 83 -572 99 -538
rect 157 -572 173 -538
rect 211 -572 227 -538
rect 353 -640 387 -578
rect -387 -674 -291 -640
rect 291 -674 387 -640
<< viali >>
rect -211 538 -173 572
rect -83 538 -45 572
rect 45 538 83 572
rect 173 538 211 572
rect -273 -488 -239 488
rect -145 -488 -111 488
rect -17 -488 17 488
rect 111 -488 145 488
rect 239 -488 273 488
rect -211 -572 -173 -538
rect -83 -572 -45 -538
rect 45 -572 83 -538
rect 173 -572 211 -538
<< metal1 >>
rect -223 572 -161 578
rect -223 538 -211 572
rect -173 538 -161 572
rect -223 532 -161 538
rect -95 572 -33 578
rect -95 538 -83 572
rect -45 538 -33 572
rect -95 532 -33 538
rect 33 572 95 578
rect 33 538 45 572
rect 83 538 95 572
rect 33 532 95 538
rect 161 572 223 578
rect 161 538 173 572
rect 211 538 223 572
rect 161 532 223 538
rect -279 488 -233 500
rect -279 -488 -273 488
rect -239 -488 -233 488
rect -279 -500 -233 -488
rect -151 488 -105 500
rect -151 -488 -145 488
rect -111 -488 -105 488
rect -151 -500 -105 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 105 488 151 500
rect 105 -488 111 488
rect 145 -488 151 488
rect 105 -500 151 -488
rect 233 488 279 500
rect 233 -488 239 488
rect 273 -488 279 488
rect 233 -500 279 -488
rect -223 -538 -161 -532
rect -223 -572 -211 -538
rect -173 -572 -161 -538
rect -223 -578 -161 -572
rect -95 -538 -33 -532
rect -95 -572 -83 -538
rect -45 -572 -33 -538
rect -95 -578 -33 -572
rect 33 -538 95 -532
rect 33 -572 45 -538
rect 83 -572 95 -538
rect 33 -578 95 -572
rect 161 -538 223 -532
rect 161 -572 173 -538
rect 211 -572 223 -538
rect 161 -578 223 -572
<< properties >>
string FIXED_BBOX -370 -657 370 657
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.0 l 0.35 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
