magic
tech sky130A
magscale 1 2
timestamp 1711565985
<< error_p >>
rect 64956 50588 65002 50600
rect 64956 50550 64962 50588
rect 64956 50538 65002 50550
rect 64956 50460 65002 50472
rect 64956 50422 64962 50460
rect 64956 50410 65002 50422
rect 64956 50332 65002 50344
rect 64956 50294 64962 50332
rect 64956 50282 65002 50294
rect 64956 50204 65002 50216
rect 64956 50166 64962 50204
rect 64956 50154 65002 50166
rect 64956 50076 65002 50088
rect 64956 50038 64962 50076
rect 64956 50026 65002 50038
rect 64956 49948 65002 49960
rect 64956 49910 64962 49948
rect 64956 49898 65002 49910
rect 64956 49820 65002 49832
rect 64956 49782 64962 49820
rect 64956 49770 65002 49782
rect 64956 49692 65002 49704
rect 64956 49654 64962 49692
rect 64956 49642 65002 49654
rect 75266 48716 75312 48728
rect 77394 48716 77440 48728
rect 77502 48716 77548 48728
rect 79630 48716 79676 48728
rect 79738 48716 79784 48728
rect 81866 48716 81912 48728
rect 75266 48678 75272 48716
rect 77394 48678 77400 48716
rect 77502 48678 77508 48716
rect 79630 48678 79636 48716
rect 79738 48678 79744 48716
rect 81866 48678 81872 48716
rect 75266 48666 75312 48678
rect 77394 48666 77440 48678
rect 77502 48666 77548 48678
rect 79630 48666 79676 48678
rect 79738 48666 79784 48678
rect 81866 48666 81912 48678
rect 77662 47158 77708 47170
rect 77770 47158 77816 47170
rect 79898 47158 79944 47170
rect 80006 47158 80052 47170
rect 82134 47158 82180 47170
rect 77662 47120 77668 47158
rect 77770 47120 77776 47158
rect 79898 47120 79904 47158
rect 80006 47120 80012 47158
rect 82134 47120 82140 47158
rect 77662 47108 77708 47120
rect 77770 47108 77816 47120
rect 79898 47108 79944 47120
rect 80006 47108 80052 47120
rect 82134 47108 82180 47120
rect 56493 45844 56539 45856
rect 57021 45844 57067 45856
rect 56493 45810 56499 45844
rect 57021 45810 57027 45844
rect 56493 45798 56539 45810
rect 57021 45798 57067 45810
rect 56493 45528 56539 45540
rect 57021 45528 57067 45540
rect 56493 45494 56499 45528
rect 57021 45494 57027 45528
rect 56493 45482 56539 45494
rect 57021 45482 57067 45494
rect 56593 45070 56639 45082
rect 56903 45070 56949 45082
rect 56593 45036 56599 45070
rect 56903 45036 56909 45070
rect 56593 45024 56639 45036
rect 56903 45024 56949 45036
rect 56593 44754 56639 44766
rect 56903 44754 56949 44766
rect 56593 44720 56599 44754
rect 56903 44720 56909 44754
rect 56593 44708 56639 44720
rect 56903 44708 56949 44720
rect 49819 41526 49865 41538
rect 50347 41526 50393 41538
rect 49819 41492 49825 41526
rect 50347 41492 50353 41526
rect 49819 41480 49865 41492
rect 50347 41480 50393 41492
rect 49819 41210 49865 41222
rect 50347 41210 50393 41222
rect 49819 41176 49825 41210
rect 50347 41176 50353 41210
rect 49819 41164 49865 41176
rect 50347 41164 50393 41176
rect 49919 40752 49965 40764
rect 50229 40752 50275 40764
rect 49919 40718 49925 40752
rect 50229 40718 50235 40752
rect 49919 40706 49965 40718
rect 50229 40706 50275 40718
rect 49919 40436 49965 40448
rect 50229 40436 50275 40448
rect 49919 40402 49925 40436
rect 50229 40402 50235 40436
rect 49919 40390 49965 40402
rect 50229 40390 50275 40402
rect 69339 31444 69401 31450
rect 69339 31410 69351 31444
rect 69339 31404 69401 31410
rect 69339 30334 69401 30340
rect 69339 30300 69351 30334
rect 69339 30294 69401 30300
rect 69339 30226 69401 30232
rect 69339 30192 69351 30226
rect 69339 30186 69401 30192
rect 53586 30011 53807 30021
rect 53840 29383 54061 30011
rect 54241 28973 54262 29779
rect 54269 29373 54516 30011
rect 54269 28945 54290 29373
rect 54670 28973 54691 29779
rect 54698 29373 54945 30011
rect 54698 28945 54719 29373
rect 55099 28973 55120 29779
rect 55127 29373 55374 30011
rect 55127 28945 55148 29373
rect 55528 28973 55549 29779
rect 55556 29373 55803 30011
rect 55556 28945 55577 29373
rect 55957 28973 55978 29779
rect 55985 29373 56232 30011
rect 55985 28945 56006 29373
rect 69339 29116 69401 29122
rect 69339 29082 69351 29116
rect 69339 29076 69401 29082
rect 69339 29008 69401 29014
rect 69339 28974 69351 29008
rect 69339 28968 69401 28974
rect 62658 28363 62692 28381
rect 62622 26904 62692 28363
rect 69339 27898 69401 27904
rect 69339 27864 69351 27898
rect 69339 27858 69401 27864
rect 69339 27790 69401 27796
rect 69339 27756 69351 27790
rect 69339 27750 69401 27756
rect 62622 26899 62693 26904
rect 62622 26863 62675 26899
rect 69339 26680 69401 26686
rect 69339 26646 69351 26680
rect 69339 26640 69401 26646
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 1000 500 44152
rect 9800 1000 10100 44152
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 200
use timer_core  timer_core_0
timestamp 1711565985
transform 1 0 45093 0 1 26552
box 0 -4258 53474 24048
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
