magic
tech sky130A
magscale 1 2
timestamp 1711842654
<< nwell >>
rect -1199 964 -823 1620
<< pwell >>
rect -1199 540 -823 964
<< nmos >>
rect -1074 628 -1044 828
rect -986 628 -956 828
<< ndiff >>
rect -1132 816 -1074 828
rect -1132 640 -1120 816
rect -1086 640 -1074 816
rect -1132 628 -1074 640
rect -1044 816 -986 828
rect -1044 639 -1032 816
rect -998 639 -986 816
rect -1044 628 -986 639
rect -956 816 -898 828
rect -956 639 -944 816
rect -910 639 -898 816
rect -956 628 -898 639
<< ndiffc >>
rect -1120 640 -1086 816
rect -1032 639 -998 816
rect -944 639 -910 816
<< psubdiff >>
rect -1163 540 -1138 574
rect -892 540 -868 574
<< nsubdiff >>
rect -1154 1550 -1130 1584
rect -892 1550 -868 1584
<< psubdiffcont >>
rect -1138 540 -892 574
<< nsubdiffcont >>
rect -1130 1550 -892 1584
<< poly >>
rect -1073 1048 -1044 1072
rect -1073 1041 -1043 1048
rect -1094 1025 -1028 1041
rect -1094 991 -1078 1025
rect -1044 991 -1028 1025
rect -1094 975 -1028 991
rect -1074 828 -1044 975
rect -985 935 -955 1072
rect -1002 919 -936 935
rect -1002 885 -986 919
rect -952 885 -936 919
rect -1002 869 -936 885
rect -986 866 -952 869
rect -986 828 -956 866
rect -1074 602 -1044 628
rect -986 602 -956 628
<< polycont >>
rect -1078 991 -1044 1025
rect -986 885 -952 919
<< locali >>
rect -1146 1550 -1130 1584
rect -892 1550 -876 1584
rect -1094 991 -1078 1025
rect -1044 991 -1028 1025
rect -1074 972 -1040 991
rect -1002 885 -986 919
rect -952 885 -936 919
rect -982 866 -948 885
rect -1120 816 -1086 832
rect -1120 624 -1086 640
rect -1032 816 -998 832
rect -944 816 -910 832
rect -1032 574 -998 639
rect -946 639 -944 816
rect -910 639 -908 816
rect -946 623 -908 639
rect -1156 540 -1138 574
rect -892 540 -876 574
<< viali >>
rect -1130 1550 -892 1584
rect -1119 1084 -1085 1460
rect -943 1084 -909 1460
rect -1078 991 -1044 1025
rect -986 885 -952 919
rect -1120 640 -1086 816
rect -944 639 -910 816
rect -1138 540 -892 574
<< metal1 >>
rect -1142 1584 -880 1590
rect -1142 1550 -1130 1584
rect -892 1550 -880 1584
rect -1142 1544 -880 1550
rect -1120 1472 -1086 1544
rect -1125 1460 -1079 1472
rect -1125 1084 -1119 1460
rect -1085 1084 -1079 1460
rect -949 1460 -903 1472
rect -949 1098 -943 1460
rect -1125 1072 -1079 1084
rect -950 1084 -943 1098
rect -909 1098 -903 1460
rect -909 1084 -877 1098
rect -950 1068 -877 1084
rect -1095 1025 -1027 1042
rect -1199 991 -1078 1025
rect -1044 991 -1027 1025
rect -1095 974 -1027 991
rect -907 1025 -877 1068
rect -907 991 -823 1025
rect -1003 919 -935 936
rect -1199 885 -986 919
rect -952 885 -935 919
rect -1003 868 -935 885
rect -907 832 -877 991
rect -1120 828 -877 832
rect -1126 816 -877 828
rect -1126 640 -1120 816
rect -1086 802 -944 816
rect -1086 640 -1080 802
rect -1126 628 -1080 640
rect -950 639 -944 802
rect -910 802 -877 816
rect -910 639 -904 802
rect -950 627 -904 639
rect -1150 574 -880 580
rect -1150 540 -1138 574
rect -892 540 -880 574
rect -1150 534 -880 540
use sky130_fd_pr__pfet_01v8_7P3MHC  sky130_fd_pr__pfet_01v8_7P3MHC_1
timestamp 1711841734
transform -1 0 -971 0 1 1236
box -141 -200 138 276
use sky130_fd_pr__pfet_01v8_7P3MHC  sky130_fd_pr__pfet_01v8_7P3MHC_2
timestamp 1711841734
transform -1 0 -1059 0 1 1236
box -141 -200 138 276
<< labels >>
flabel metal1 -1199 991 -1165 1025 3 FreeSans 160 0 0 0 IN_A
port 0 e default input
flabel metal1 -1199 885 -1165 919 3 FreeSans 160 0 0 0 IN_B
port 1 e default input
flabel metal1 -857 991 -823 1025 7 FreeSans 160 0 0 0 OUT
port 2 w default output
flabel metal1 -1130 1550 -892 1584 0 FreeSans 320 0 0 0 vdd
port 3 nsew default bidirectional
flabel metal1 -1138 540 -892 574 0 FreeSans 320 0 0 0 vss
port 4 nsew default bidirectional
<< end >>
