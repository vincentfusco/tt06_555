magic
tech sky130A
magscale 1 2
timestamp 1710860902
<< pwell >>
rect -296 -2319 296 2319
<< nmos >>
rect -100 109 100 2109
rect -100 -2109 100 -109
<< ndiff >>
rect -158 2097 -100 2109
rect -158 121 -146 2097
rect -112 121 -100 2097
rect -158 109 -100 121
rect 100 2097 158 2109
rect 100 121 112 2097
rect 146 121 158 2097
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -2097 -146 -121
rect -112 -2097 -100 -121
rect -158 -2109 -100 -2097
rect 100 -121 158 -109
rect 100 -2097 112 -121
rect 146 -2097 158 -121
rect 100 -2109 158 -2097
<< ndiffc >>
rect -146 121 -112 2097
rect 112 121 146 2097
rect -146 -2097 -112 -121
rect 112 -2097 146 -121
<< psubdiff >>
rect -260 2249 -164 2283
rect 164 2249 260 2283
rect -260 2187 -226 2249
rect 226 2187 260 2249
rect -260 -2249 -226 -2187
rect 226 -2249 260 -2187
rect -260 -2283 -164 -2249
rect 164 -2283 260 -2249
<< psubdiffcont >>
rect -164 2249 164 2283
rect -260 -2187 -226 2187
rect 226 -2187 260 2187
rect -164 -2283 164 -2249
<< poly >>
rect -100 2181 100 2197
rect -100 2147 -84 2181
rect 84 2147 100 2181
rect -100 2109 100 2147
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -2147 100 -2109
rect -100 -2181 -84 -2147
rect 84 -2181 100 -2147
rect -100 -2197 100 -2181
<< polycont >>
rect -84 2147 84 2181
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -2181 84 -2147
<< locali >>
rect -260 2249 -164 2283
rect 164 2249 260 2283
rect -260 2187 -226 2249
rect 226 2187 260 2249
rect -100 2147 -84 2181
rect 84 2147 100 2181
rect -146 2097 -112 2113
rect -146 105 -112 121
rect 112 2097 146 2113
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -2113 -112 -2097
rect 112 -121 146 -105
rect 112 -2113 146 -2097
rect -100 -2181 -84 -2147
rect 84 -2181 100 -2147
rect -260 -2249 -226 -2187
rect 226 -2249 260 -2187
rect -260 -2283 -164 -2249
rect 164 -2283 260 -2249
<< viali >>
rect -84 2147 84 2181
rect -146 121 -112 2097
rect 112 121 146 2097
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -2097 -112 -121
rect 112 -2097 146 -121
rect -84 -2181 84 -2147
<< metal1 >>
rect -96 2181 96 2187
rect -96 2147 -84 2181
rect 84 2147 96 2181
rect -96 2141 96 2147
rect -152 2097 -106 2109
rect -152 121 -146 2097
rect -112 121 -106 2097
rect -152 109 -106 121
rect 106 2097 152 2109
rect 106 121 112 2097
rect 146 121 152 2097
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -2097 -146 -121
rect -112 -2097 -106 -121
rect -152 -2109 -106 -2097
rect 106 -121 152 -109
rect 106 -2097 112 -121
rect 146 -2097 152 -121
rect 106 -2109 152 -2097
rect -96 -2147 96 -2141
rect -96 -2181 -84 -2147
rect 84 -2181 96 -2147
rect -96 -2187 96 -2181
<< properties >>
string FIXED_BBOX -243 -2266 243 2266
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
