magic
tech sky130A
magscale 1 2
timestamp 1711041017
<< error_p >>
rect -31 2399 31 2405
rect -31 2365 -19 2399
rect -31 2359 31 2365
rect -31 1289 31 1295
rect -31 1255 -19 1289
rect -31 1249 31 1255
rect -31 1181 31 1187
rect -31 1147 -19 1181
rect -31 1141 31 1147
rect -31 71 31 77
rect -31 37 -19 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect -31 -77 31 -71
rect -31 -1147 31 -1141
rect -31 -1181 -19 -1147
rect -31 -1187 31 -1181
rect -31 -1255 31 -1249
rect -31 -1289 -19 -1255
rect -31 -1295 31 -1289
rect -31 -2365 31 -2359
rect -31 -2399 -19 -2365
rect -31 -2405 31 -2399
<< pwell >>
rect -231 -2537 2431 2537
<< nmoslvt >>
rect -35 1327 35 2327
rect -35 109 35 1109
rect -35 -1109 35 -109
rect -35 -2327 35 -1327
<< ndiff >>
rect -93 2315 -35 2327
rect -93 1339 -81 2315
rect -47 1339 -35 2315
rect -93 1327 -35 1339
rect 35 2315 93 2327
rect 35 1339 47 2315
rect 81 1339 93 2315
rect 35 1327 93 1339
rect -93 1097 -35 1109
rect -93 121 -81 1097
rect -47 121 -35 1097
rect -93 109 -35 121
rect 35 1097 93 1109
rect 35 121 47 1097
rect 81 121 93 1097
rect 35 109 93 121
rect -93 -121 -35 -109
rect -93 -1097 -81 -121
rect -47 -1097 -35 -121
rect -93 -1109 -35 -1097
rect 35 -121 93 -109
rect 35 -1097 47 -121
rect 81 -1097 93 -121
rect 35 -1109 93 -1097
rect -93 -1339 -35 -1327
rect -93 -2315 -81 -1339
rect -47 -2315 -35 -1339
rect -93 -2327 -35 -2315
rect 35 -1339 93 -1327
rect 35 -2315 47 -1339
rect 81 -2315 93 -1339
rect 35 -2327 93 -2315
<< ndiffc >>
rect -81 1339 -47 2315
rect 47 1339 81 2315
rect -81 121 -47 1097
rect 47 121 81 1097
rect -81 -1097 -47 -121
rect 47 -1097 81 -121
rect -81 -2315 -47 -1339
rect 47 -2315 81 -1339
<< psubdiff >>
rect -195 2467 -99 2501
rect 99 2467 2395 2501
rect -195 2405 -161 2467
rect 2361 2405 2395 2467
rect -195 -2467 -161 -2405
rect 2361 -2467 2395 -2405
rect -195 -2501 -99 -2467
rect 99 -2501 2395 -2467
<< psubdiffcont >>
rect -99 2467 99 2501
rect -195 -2405 -161 2405
rect 2361 -2405 2395 2405
rect -99 -2501 99 -2467
<< poly >>
rect -35 2399 35 2415
rect -35 2365 -19 2399
rect 19 2365 35 2399
rect -35 2327 35 2365
rect -35 1289 35 1327
rect -35 1255 -19 1289
rect 19 1255 35 1289
rect -35 1239 35 1255
rect -35 1181 35 1197
rect -35 1147 -19 1181
rect 19 1147 35 1181
rect -35 1109 35 1147
rect -35 71 35 109
rect -35 37 -19 71
rect 19 37 35 71
rect -35 21 35 37
rect -35 -37 35 -21
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect -35 -109 35 -71
rect -35 -1147 35 -1109
rect -35 -1181 -19 -1147
rect 19 -1181 35 -1147
rect -35 -1197 35 -1181
rect -35 -1255 35 -1239
rect -35 -1289 -19 -1255
rect 19 -1289 35 -1255
rect -35 -1327 35 -1289
rect -35 -2365 35 -2327
rect -35 -2399 -19 -2365
rect 19 -2399 35 -2365
rect -35 -2415 35 -2399
<< polycont >>
rect -19 2365 19 2399
rect -19 1255 19 1289
rect -19 1147 19 1181
rect -19 37 19 71
rect -19 -71 19 -37
rect -19 -1181 19 -1147
rect -19 -1289 19 -1255
rect -19 -2399 19 -2365
<< locali >>
rect -195 2467 -99 2501
rect 99 2467 2395 2501
rect -195 2405 -161 2467
rect 2361 2405 2395 2467
rect -35 2365 -19 2399
rect 19 2365 35 2399
rect -81 2315 -47 2331
rect -81 1323 -47 1339
rect 47 2315 81 2331
rect 47 1323 81 1339
rect -35 1255 -19 1289
rect 19 1255 35 1289
rect -35 1147 -19 1181
rect 19 1147 35 1181
rect -81 1097 -47 1113
rect -81 105 -47 121
rect 47 1097 81 1113
rect 47 105 81 121
rect -35 37 -19 71
rect 19 37 35 71
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect -81 -121 -47 -105
rect -81 -1113 -47 -1097
rect 47 -121 81 -105
rect 47 -1113 81 -1097
rect -35 -1181 -19 -1147
rect 19 -1181 35 -1147
rect -35 -1289 -19 -1255
rect 19 -1289 35 -1255
rect -81 -1339 -47 -1323
rect -81 -2331 -47 -2315
rect 47 -1339 81 -1323
rect 47 -2331 81 -2315
rect -35 -2399 -19 -2365
rect 19 -2399 35 -2365
rect -195 -2467 -161 -2405
rect 2361 -2467 2395 -2405
rect -195 -2501 -99 -2467
rect 99 -2501 2395 -2467
<< viali >>
rect -19 2365 19 2399
rect -81 1339 -47 2315
rect 47 1339 81 2315
rect -19 1255 19 1289
rect -19 1147 19 1181
rect -81 121 -47 1097
rect 47 121 81 1097
rect -19 37 19 71
rect -19 -71 19 -37
rect -81 -1097 -47 -121
rect 47 -1097 81 -121
rect -19 -1181 19 -1147
rect -19 -1289 19 -1255
rect -81 -2315 -47 -1339
rect 47 -2315 81 -1339
rect -19 -2399 19 -2365
<< metal1 >>
rect -31 2399 31 2405
rect -31 2365 -19 2399
rect 19 2365 31 2399
rect -31 2359 31 2365
rect -87 2315 -41 2327
rect -87 1339 -81 2315
rect -47 1339 -41 2315
rect -87 1327 -41 1339
rect 41 2315 87 2327
rect 41 1339 47 2315
rect 81 1339 87 2315
rect 41 1327 87 1339
rect -31 1289 31 1295
rect -31 1255 -19 1289
rect 19 1255 31 1289
rect -31 1249 31 1255
rect -31 1181 31 1187
rect -31 1147 -19 1181
rect 19 1147 31 1181
rect -31 1141 31 1147
rect -87 1097 -41 1109
rect -87 121 -81 1097
rect -47 121 -41 1097
rect -87 109 -41 121
rect 41 1097 87 1109
rect 41 121 47 1097
rect 81 121 87 1097
rect 41 109 87 121
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect -87 -121 -41 -109
rect -87 -1097 -81 -121
rect -47 -1097 -41 -121
rect -87 -1109 -41 -1097
rect 41 -121 87 -109
rect 41 -1097 47 -121
rect 81 -1097 87 -121
rect 41 -1109 87 -1097
rect -31 -1147 31 -1141
rect -31 -1181 -19 -1147
rect 19 -1181 31 -1147
rect -31 -1187 31 -1181
rect -31 -1255 31 -1249
rect -31 -1289 -19 -1255
rect 19 -1289 31 -1255
rect -31 -1295 31 -1289
rect -87 -1339 -41 -1327
rect -87 -2315 -81 -1339
rect -47 -2315 -41 -1339
rect -87 -2327 -41 -2315
rect 41 -1339 87 -1327
rect 41 -2315 47 -1339
rect 81 -2315 87 -1339
rect 41 -2327 87 -2315
rect -31 -2365 31 -2359
rect -31 -2399 -19 -2365
rect 19 -2399 31 -2365
rect -31 -2405 31 -2399
<< properties >>
string FIXED_BBOX -178 -2484 178 2484
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.0 l 0.35 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
