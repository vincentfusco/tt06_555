magic
tech sky130A
magscale 1 2
timestamp 1711045747
<< error_p >>
rect 2655 5236 2701 5248
rect 3183 5236 3229 5248
rect 2655 5202 2661 5236
rect 3183 5202 3189 5236
rect 2655 5190 2701 5202
rect 3183 5190 3229 5202
rect 2655 4920 2701 4932
rect 3183 4920 3229 4932
rect 2655 4886 2661 4920
rect 3183 4886 3189 4920
rect 2655 4874 2701 4886
rect 3183 4874 3229 4886
rect 2755 4462 2801 4474
rect 3065 4462 3111 4474
rect 2755 4428 2761 4462
rect 3065 4428 3071 4462
rect 2755 4416 2801 4428
rect 3065 4416 3111 4428
rect 2755 4146 2801 4158
rect 3065 4146 3111 4158
rect 2755 4112 2761 4146
rect 3065 4112 3071 4146
rect 2755 4100 2801 4112
rect 3065 4100 3111 4112
rect -4019 918 -3973 930
rect -3491 918 -3445 930
rect -4019 884 -4013 918
rect -3491 884 -3485 918
rect -4019 872 -3973 884
rect -3491 872 -3445 884
rect -4019 602 -3973 614
rect -3491 602 -3445 614
rect -4019 568 -4013 602
rect -3491 568 -3485 602
rect -4019 556 -3973 568
rect -3491 556 -3445 568
rect -3919 144 -3873 156
rect -3609 144 -3563 156
rect -3919 110 -3913 144
rect -3609 110 -3603 144
rect -3919 98 -3873 110
rect -3609 98 -3563 110
rect -3919 -172 -3873 -160
rect -3609 -172 -3563 -160
rect -3919 -206 -3913 -172
rect -3609 -206 -3603 -172
rect -3919 -218 -3873 -206
rect -3609 -218 -3563 -206
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use nor  X_NOR_R
timestamp 1711045747
transform 1 0 1853 0 1 4138
box 364 -1040 1850 1568
use nor  X_NOR_S1
timestamp 1711045747
transform 1 0 -4821 0 1 -180
box 364 -1040 1850 1568
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 IN_S
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 OUT_Q_B
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 IN_R
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 OUT_Q
port 5 nsew
<< end >>
