magic
tech sky130A
magscale 1 2
timestamp 1711736161
<< error_p >>
rect -159 1072 -97 1078
rect -31 1072 31 1078
rect 97 1072 159 1078
rect -159 1038 -147 1072
rect -31 1038 -19 1072
rect 97 1038 109 1072
rect -159 1032 -97 1038
rect -31 1032 31 1038
rect 97 1032 159 1038
rect -159 -1038 -97 -1032
rect -31 -1038 31 -1032
rect 97 -1038 159 -1032
rect -159 -1072 -147 -1038
rect -31 -1072 -19 -1038
rect 97 -1072 109 -1038
rect -159 -1078 -97 -1072
rect -31 -1078 31 -1072
rect 97 -1078 159 -1072
<< pwell >>
rect -359 -1210 359 1210
<< nmoslvt >>
rect -163 -1000 -93 1000
rect -35 -1000 35 1000
rect 93 -1000 163 1000
<< ndiff >>
rect -221 988 -163 1000
rect -221 -988 -209 988
rect -175 -988 -163 988
rect -221 -1000 -163 -988
rect -93 988 -35 1000
rect -93 -988 -81 988
rect -47 -988 -35 988
rect -93 -1000 -35 -988
rect 35 988 93 1000
rect 35 -988 47 988
rect 81 -988 93 988
rect 35 -1000 93 -988
rect 163 988 221 1000
rect 163 -988 175 988
rect 209 -988 221 988
rect 163 -1000 221 -988
<< ndiffc >>
rect -209 -988 -175 988
rect -81 -988 -47 988
rect 47 -988 81 988
rect 175 -988 209 988
<< psubdiff >>
rect -323 1140 -227 1174
rect 227 1140 323 1174
rect -323 1078 -289 1140
rect 289 1078 323 1140
rect -323 -1140 -289 -1078
rect 289 -1140 323 -1078
rect -323 -1174 -227 -1140
rect 227 -1174 323 -1140
<< psubdiffcont >>
rect -227 1140 227 1174
rect -323 -1078 -289 1078
rect 289 -1078 323 1078
rect -227 -1174 227 -1140
<< poly >>
rect -163 1072 -93 1088
rect -163 1038 -147 1072
rect -109 1038 -93 1072
rect -163 1000 -93 1038
rect -35 1072 35 1088
rect -35 1038 -19 1072
rect 19 1038 35 1072
rect -35 1000 35 1038
rect 93 1072 163 1088
rect 93 1038 109 1072
rect 147 1038 163 1072
rect 93 1000 163 1038
rect -163 -1038 -93 -1000
rect -163 -1072 -147 -1038
rect -109 -1072 -93 -1038
rect -163 -1088 -93 -1072
rect -35 -1038 35 -1000
rect -35 -1072 -19 -1038
rect 19 -1072 35 -1038
rect -35 -1088 35 -1072
rect 93 -1038 163 -1000
rect 93 -1072 109 -1038
rect 147 -1072 163 -1038
rect 93 -1088 163 -1072
<< polycont >>
rect -147 1038 -109 1072
rect -19 1038 19 1072
rect 109 1038 147 1072
rect -147 -1072 -109 -1038
rect -19 -1072 19 -1038
rect 109 -1072 147 -1038
<< locali >>
rect -323 1140 -227 1174
rect 227 1140 323 1174
rect -323 1078 -289 1140
rect 289 1078 323 1140
rect -163 1038 -147 1072
rect -109 1038 -93 1072
rect -35 1038 -19 1072
rect 19 1038 35 1072
rect 93 1038 109 1072
rect 147 1038 163 1072
rect -209 988 -175 1004
rect -209 -1004 -175 -988
rect -81 988 -47 1004
rect -81 -1004 -47 -988
rect 47 988 81 1004
rect 47 -1004 81 -988
rect 175 988 209 1004
rect 175 -1004 209 -988
rect -163 -1072 -147 -1038
rect -109 -1072 -93 -1038
rect -35 -1072 -19 -1038
rect 19 -1072 35 -1038
rect 93 -1072 109 -1038
rect 147 -1072 163 -1038
rect -323 -1140 -289 -1078
rect 289 -1140 323 -1078
rect -323 -1174 -227 -1140
rect 227 -1174 323 -1140
<< viali >>
rect -147 1038 -109 1072
rect -19 1038 19 1072
rect 109 1038 147 1072
rect -209 -988 -175 988
rect -81 -988 -47 988
rect 47 -988 81 988
rect 175 -988 209 988
rect -147 -1072 -109 -1038
rect -19 -1072 19 -1038
rect 109 -1072 147 -1038
<< metal1 >>
rect -159 1072 -97 1078
rect -159 1038 -147 1072
rect -109 1038 -97 1072
rect -159 1032 -97 1038
rect -31 1072 31 1078
rect -31 1038 -19 1072
rect 19 1038 31 1072
rect -31 1032 31 1038
rect 97 1072 159 1078
rect 97 1038 109 1072
rect 147 1038 159 1072
rect 97 1032 159 1038
rect -215 988 -169 1000
rect -215 -988 -209 988
rect -175 -988 -169 988
rect -215 -1000 -169 -988
rect -87 988 -41 1000
rect -87 -988 -81 988
rect -47 -988 -41 988
rect -87 -1000 -41 -988
rect 41 988 87 1000
rect 41 -988 47 988
rect 81 -988 87 988
rect 41 -1000 87 -988
rect 169 988 215 1000
rect 169 -988 175 988
rect 209 -988 215 988
rect 169 -1000 215 -988
rect -159 -1038 -97 -1032
rect -159 -1072 -147 -1038
rect -109 -1072 -97 -1038
rect -159 -1078 -97 -1072
rect -31 -1038 31 -1032
rect -31 -1072 -19 -1038
rect 19 -1072 31 -1038
rect -31 -1078 31 -1072
rect 97 -1038 159 -1032
rect 97 -1072 109 -1038
rect 147 -1072 159 -1038
rect 97 -1078 159 -1072
<< properties >>
string FIXED_BBOX -306 -1157 306 1157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 10 l 0.35 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
