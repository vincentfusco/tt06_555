magic
tech sky130A
magscale 1 2
timestamp 1710860643
<< nwell >>
rect -296 -2337 296 2337
<< pmos >>
rect -100 118 100 2118
rect -100 -2118 100 -118
<< pdiff >>
rect -158 2106 -100 2118
rect -158 130 -146 2106
rect -112 130 -100 2106
rect -158 118 -100 130
rect 100 2106 158 2118
rect 100 130 112 2106
rect 146 130 158 2106
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -2106 -146 -130
rect -112 -2106 -100 -130
rect -158 -2118 -100 -2106
rect 100 -130 158 -118
rect 100 -2106 112 -130
rect 146 -2106 158 -130
rect 100 -2118 158 -2106
<< pdiffc >>
rect -146 130 -112 2106
rect 112 130 146 2106
rect -146 -2106 -112 -130
rect 112 -2106 146 -130
<< nsubdiff >>
rect -260 2267 -164 2301
rect 164 2267 260 2301
rect -260 2205 -226 2267
rect 226 2205 260 2267
rect -260 -2267 -226 -2205
rect 226 -2267 260 -2205
rect -260 -2301 -164 -2267
rect 164 -2301 260 -2267
<< nsubdiffcont >>
rect -164 2267 164 2301
rect -260 -2205 -226 2205
rect 226 -2205 260 2205
rect -164 -2301 164 -2267
<< poly >>
rect -100 2199 100 2215
rect -100 2165 -84 2199
rect 84 2165 100 2199
rect -100 2118 100 2165
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -2165 100 -2118
rect -100 -2199 -84 -2165
rect 84 -2199 100 -2165
rect -100 -2215 100 -2199
<< polycont >>
rect -84 2165 84 2199
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -2199 84 -2165
<< locali >>
rect -260 2267 -164 2301
rect 164 2267 260 2301
rect -260 2205 -226 2267
rect 226 2205 260 2267
rect -100 2165 -84 2199
rect 84 2165 100 2199
rect -146 2106 -112 2122
rect -146 114 -112 130
rect 112 2106 146 2122
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -2122 -112 -2106
rect 112 -130 146 -114
rect 112 -2122 146 -2106
rect -100 -2199 -84 -2165
rect 84 -2199 100 -2165
rect -260 -2267 -226 -2205
rect 226 -2267 260 -2205
rect -260 -2301 -164 -2267
rect 164 -2301 260 -2267
<< viali >>
rect -84 2165 84 2199
rect -146 130 -112 2106
rect 112 130 146 2106
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -2106 -112 -130
rect 112 -2106 146 -130
rect -84 -2199 84 -2165
<< metal1 >>
rect -96 2199 96 2205
rect -96 2165 -84 2199
rect 84 2165 96 2199
rect -96 2159 96 2165
rect -152 2106 -106 2118
rect -152 130 -146 2106
rect -112 130 -106 2106
rect -152 118 -106 130
rect 106 2106 152 2118
rect 106 130 112 2106
rect 146 130 152 2106
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -2106 -146 -130
rect -112 -2106 -106 -130
rect -152 -2118 -106 -2106
rect 106 -130 152 -118
rect 106 -2106 112 -130
rect 146 -2106 152 -130
rect 106 -2118 152 -2106
rect -96 -2165 96 -2159
rect -96 -2199 -84 -2165
rect 84 -2199 96 -2165
rect -96 -2205 96 -2199
<< properties >>
string FIXED_BBOX -243 -2284 243 2284
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
