magic
tech sky130A
magscale 1 2
timestamp 1711041017
<< nmoslvt >>
rect -227 -500 -157 500
rect -99 -500 -29 500
rect 29 -500 99 500
rect 157 -500 227 500
<< ndiff >>
rect -285 488 -227 500
rect -285 -488 -273 488
rect -239 -488 -227 488
rect -285 -500 -227 -488
rect -157 488 -99 500
rect -157 -488 -145 488
rect -111 -488 -99 488
rect -157 -500 -99 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 99 488 157 500
rect 99 -488 111 488
rect 145 -488 157 488
rect 99 -500 157 -488
rect 227 488 285 500
rect 227 -488 239 488
rect 273 -488 285 488
rect 227 -500 285 -488
<< ndiffc >>
rect -273 -488 -239 488
rect -145 -488 -111 488
rect -17 -488 17 488
rect 111 -488 145 488
rect 239 -488 273 488
<< poly >>
rect -227 500 -157 526
rect -99 500 -29 526
rect 29 500 99 526
rect 157 500 227 526
rect -227 -526 -157 -500
rect -99 -526 -29 -500
rect 29 -526 99 -500
rect 157 -526 227 -500
<< locali >>
rect -273 488 -239 504
rect -273 -504 -239 -488
rect -145 488 -111 504
rect -145 -504 -111 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 111 488 145 504
rect 111 -504 145 -488
rect 239 488 273 504
rect 239 -504 273 -488
<< viali >>
rect -273 -488 -239 488
rect -145 -488 -111 488
rect -17 -488 17 488
rect 111 -488 145 488
rect 239 -488 273 488
<< metal1 >>
rect -279 488 -233 500
rect -279 -488 -273 488
rect -239 -488 -233 488
rect -279 -500 -233 -488
rect -151 488 -105 500
rect -151 -488 -145 488
rect -111 -488 -105 488
rect -151 -500 -105 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 105 488 151 500
rect 105 -488 111 488
rect 145 -488 151 488
rect 105 -500 151 -488
rect 233 488 279 500
rect 233 -488 239 488
rect 273 -488 279 488
rect 233 -500 279 -488
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.0 l 0.35 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
