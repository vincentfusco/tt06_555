* NGSPICE file created from tt_um_vaf_555_timer.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_BXYDM4 a_15_n131# a_n15_n157# a_n73_n131# VSUBS
X0 a_15_n131# a_n15_n157# a_n73_n131# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n73_n131# a_15_n131# 0.166179f
C1 a_n15_n157# a_15_n131# 0.013387f
C2 a_n15_n157# a_n73_n131# 0.005542f
C3 a_15_n131# VSUBS 0.116709f
C4 a_n73_n131# VSUBS 0.118252f
C5 a_n15_n157# VSUBS 0.066041f
.ends

.subckt sky130_fd_pr__pfet_01v8_7PK3FC a_n73_n64# a_n33_n161# m1_n141_190# a_15_n64#
+ w_n141_n178# VSUBS
X0 a_15_n64# a_n33_n161# a_n73_n64# w_n141_n178# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_15_n64# m1_n141_190# 0.020547f
C1 a_n73_n64# m1_n141_190# 0.020547f
C2 a_n33_n161# m1_n141_190# 0.009013f
C3 a_n73_n64# a_15_n64# 0.162113f
C4 a_n33_n161# a_15_n64# 0.017761f
C5 w_n141_n178# m1_n141_190# 0.046696f
C6 w_n141_n178# a_15_n64# 0.021345f
C7 a_n33_n161# a_n73_n64# 0.017761f
C8 w_n141_n178# a_n73_n64# 0.021345f
C9 w_n141_n178# a_n33_n161# 0.084351f
C10 m1_n141_190# VSUBS 0.083142f
C11 a_15_n64# VSUBS 0.089867f
C12 a_n73_n64# VSUBS 0.089867f
C13 a_n33_n161# VSUBS 0.130601f
C14 w_n141_n178# VSUBS 0.464632f
.ends

.subckt inv vout vss vdd vin
XXMn vout vin vss vss sky130_fd_pr__nfet_01v8_BXYDM4
Xsky130_fd_pr__pfet_01v8_7PK3FC_0 vdd vin vdd vout vdd vss sky130_fd_pr__pfet_01v8_7PK3FC
C0 vout vdd 0.069903f
C1 vss vdd 0.005257f
C2 vin vdd 0.07994f
C3 vss vout -0.06331f
C4 vin vout 0.13222f
C5 vin vss 0.011685f
C6 vdd 0 0.815242f
C7 vout 0 0.442391f
C8 vss 0 0.026556f
C9 vin 0 0.446699f
.ends

.subckt sky130_fd_pr__pfet_01v8_7P3MHC a_n16_n190# w_n141_n200# a_n74_n164# a_14_n164#
+ VSUBS
X0 a_14_n164# a_n16_n190# a_n74_n164# w_n141_n200# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_14_n164# a_n74_n164# 0.127297f
C1 w_n141_n200# a_n74_n164# 0.002485f
C2 a_n16_n190# a_n74_n164# 0.001584f
C3 w_n141_n200# a_14_n164# 0.002471f
C4 a_n16_n190# a_14_n164# 0.001584f
C5 a_n16_n190# w_n141_n200# 0.022362f
C6 a_14_n164# VSUBS 0.104203f
C7 a_n74_n164# VSUBS 0.104189f
C8 a_n16_n190# VSUBS 0.04368f
C9 w_n141_n200# VSUBS 0.398412f
.ends

.subckt nor IN_A IN_B OUT vdd vss sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
Xsky130_fd_pr__pfet_01v8_7P3MHC_1 IN_B vdd OUT sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ vss sky130_fd_pr__pfet_01v8_7P3MHC
Xsky130_fd_pr__pfet_01v8_7P3MHC_2 IN_A vdd sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ vdd vss sky130_fd_pr__pfet_01v8_7P3MHC
X0 OUT IN_B vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X1 vss IN_A OUT vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
C0 IN_A OUT 0.042579f
C1 sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# OUT 0.02361f
C2 vdd OUT 0.166932f
C3 IN_B OUT 0.176005f
C4 sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# IN_A 0.005339f
C5 vdd IN_A 0.117603f
C6 vdd sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 0.037594f
C7 IN_B IN_A 0.172705f
C8 IN_B sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 0.005333f
C9 IN_B vdd 0.058945f
C10 IN_A vss 0.194746f
C11 sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# vss 0.022957f
C12 OUT vss 0.689203f
C13 IN_B vss 0.229565f
C14 vdd vss 1.048658f
.ends

.subckt nand IN_A IN_B OUT vdd vss drain_mna
Xsky130_fd_pr__pfet_01v8_7P3MHC_1 IN_B vdd OUT vdd vss sky130_fd_pr__pfet_01v8_7P3MHC
Xsky130_fd_pr__pfet_01v8_7P3MHC_2 IN_A vdd vdd OUT vss sky130_fd_pr__pfet_01v8_7P3MHC
X0 OUT IN_B drain_mna vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X1 drain_mna IN_A vss vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
C0 OUT vdd 0.190223f
C1 drain_mna vdd 0.003922f
C2 IN_B vdd 0.05155f
C3 IN_A vdd 0.070703f
C4 drain_mna OUT 0.080424f
C5 IN_B OUT 0.112665f
C6 IN_A OUT 0.080949f
C7 IN_B drain_mna 0.011696f
C8 IN_A drain_mna 0.001675f
C9 IN_A IN_B 0.176887f
C10 drain_mna vss 0.108169f
C11 IN_A vss 0.207303f
C12 OUT vss 0.589588f
C13 IN_B vss 0.265243f
C14 vdd vss 0.92595f
.ends

.subckt sr_latch_rb IN_S IN_R IN_R_N OUT_Q vdd X_NOR_TOP/OUT X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ inv_0/vout nand_0/drain_mna vss nand_0/OUT X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
Xinv_0 inv_0/vout vss vdd IN_R inv
XX_NOR_TOP OUT_Q IN_S X_NOR_TOP/OUT vdd vss X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ nor
XX_NOR_BOTTOM X_NOR_TOP/OUT nand_0/OUT OUT_Q vdd vss X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ nor
Xnand_0 inv_0/vout IN_R_N nand_0/OUT vdd vss nand_0/drain_mna nand
C0 inv_0/vout nand_0/drain_mna 1.37e-19
C1 X_NOR_TOP/OUT X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 3.49e-20
C2 OUT_Q nand_0/drain_mna 4.91e-21
C3 vss IN_R_N 0.119198f
C4 IN_S IN_R_N 0.100958f
C5 X_NOR_TOP/OUT IN_R 7.13e-20
C6 inv_0/vout IN_R_N 0.101216f
C7 nand_0/OUT IN_R 0.006121f
C8 vdd IN_R 0.009435f
C9 OUT_Q IN_R_N 0.021916f
C10 X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# IN_R 6.23e-20
C11 IN_S X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 0.001116f
C12 vss IN_R -2.29e-19
C13 IN_S IN_R 0.137576f
C14 inv_0/vout IN_R 0.012448f
C15 OUT_Q X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 0.006615f
C16 IN_R_N nand_0/drain_mna 0.004493f
C17 OUT_Q IN_R 4.08e-20
C18 IN_R nand_0/drain_mna 5.17e-21
C19 IN_R IN_R_N 0.048793f
C20 IN_R X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 2.57e-20
C21 nand_0/OUT X_NOR_TOP/OUT 0.276403f
C22 vdd X_NOR_TOP/OUT 0.175916f
C23 vdd nand_0/OUT 0.16551f
C24 X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# nand_0/OUT 5.92e-20
C25 vss X_NOR_TOP/OUT 0.041485f
C26 IN_S X_NOR_TOP/OUT 0.024837f
C27 X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# vdd 2.81e-20
C28 vss nand_0/OUT 0.032732f
C29 inv_0/vout X_NOR_TOP/OUT 1.19e-19
C30 vss vdd 1.96e-19
C31 IN_S nand_0/OUT 0.349702f
C32 inv_0/vout nand_0/OUT 0.156863f
C33 IN_S vdd 0.188524f
C34 inv_0/vout vdd 0.041062f
C35 OUT_Q X_NOR_TOP/OUT 0.295691f
C36 IN_S X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 0.00251f
C37 OUT_Q nand_0/OUT 0.111763f
C38 OUT_Q vdd 0.061303f
C39 IN_S vss 0.004506f
C40 inv_0/vout vss 0.090793f
C41 OUT_Q X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 0.007086f
C42 inv_0/vout IN_S 0.194534f
C43 X_NOR_TOP/OUT nand_0/drain_mna 1.73e-19
C44 OUT_Q vss 0.001965f
C45 OUT_Q IN_S 0.096978f
C46 nand_0/OUT nand_0/drain_mna 1.91e-19
C47 OUT_Q inv_0/vout 0.003946f
C48 X_NOR_TOP/OUT IN_R_N 0.007502f
C49 vss nand_0/drain_mna 7.25e-20
C50 nand_0/OUT IN_R_N 0.01683f
C51 IN_S nand_0/drain_mna 0.003085f
C52 vdd IN_R_N 0.011685f
C53 nand_0/drain_mna 0 0.108169f
C54 nand_0/OUT 0 0.524253f
C55 IN_R_N 0 0.369798f
C56 X_NOR_TOP/OUT 0 0.629748f
C57 X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 0 0.020446f
C58 OUT_Q 0 0.835481f
C59 X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 0 0.020446f
C60 IN_S 0 0.389263f
C61 vdd 0 3.455888f
C62 inv_0/vout 0 0.382539f
C63 vss 0 -0.801757f
C64 IN_R 0 0.311523f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_MMMA4V a_n260_n698# a_100_n500# a_n158_n500# a_n100_n588#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n260_n698# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
C0 a_100_n500# a_n158_n500# 0.273876f
C1 a_n100_n588# a_n158_n500# 0.112293f
C2 a_100_n500# a_n100_n588# 0.112293f
C3 a_100_n500# a_n260_n698# 0.590504f
C4 a_n158_n500# a_n260_n698# 0.590504f
C5 a_n100_n588# a_n260_n698# 0.718303f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_5VNMZ8 a_n100_n897# a_100_n800# w_n296_n1019#
+ a_n158_n800# VSUBS
X0 a_100_n800# a_n100_n897# a_n158_n800# w_n296_n1019# sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
C0 a_n158_n800# a_n100_n897# 0.176406f
C1 a_100_n800# a_n100_n897# 0.176406f
C2 a_n158_n800# a_100_n800# 0.437576f
C3 w_n296_n1019# a_n100_n897# 0.434431f
C4 a_n158_n800# w_n296_n1019# 0.512046f
C5 w_n296_n1019# a_100_n800# 0.512046f
C6 a_100_n800# VSUBS 0.413693f
C7 a_n158_n800# VSUBS 0.413693f
C8 a_n100_n897# VSUBS 0.364183f
C9 w_n296_n1019# VSUBS 4.82082f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AHMAL2 a_n260_n574# a_100_n400# a_n158_n400# a_n100_n488#
X0 a_100_n400# a_n100_n488# a_n158_n400# a_n260_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
C0 a_100_n400# a_n158_n400# 0.219309f
C1 a_n100_n488# a_n158_n400# 0.090922f
C2 a_100_n400# a_n100_n488# 0.090922f
C3 a_100_n400# a_n260_n574# 0.480566f
C4 a_n158_n400# a_n260_n574# 0.480566f
C5 a_n100_n488# a_n260_n574# 0.74751f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_GUWLND a_n158_n1000# a_n100_n1097# w_n296_n1219#
+ a_100_n1000# VSUBS
X0 a_100_n1000# a_n100_n1097# a_n158_n1000# w_n296_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
C0 a_n158_n1000# a_n100_n1097# 0.219148f
C1 a_100_n1000# a_n100_n1097# 0.219148f
C2 a_n158_n1000# a_100_n1000# 0.54671f
C3 w_n296_n1219# a_n100_n1097# 0.434431f
C4 a_n158_n1000# w_n296_n1219# 0.633996f
C5 w_n296_n1219# a_100_n1000# 0.633996f
C6 a_100_n1000# VSUBS 0.514548f
C7 a_n158_n1000# VSUBS 0.514548f
C8 a_n100_n1097# VSUBS 0.364183f
C9 w_n296_n1219# VSUBS 5.72384f
.ends

.subckt comp_p vinp vinn vbias_p vdd latch_left tail out_left vout latch_right vss
XXMn_cs_left vss latch_right vss latch_left sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMp_out out_left vdd vdd vout vss sky130_fd_pr__pfet_01v8_lvt_5VNMZ8
XXMn_diode_left1 vss latch_left vss latch_left sky130_fd_pr__nfet_01v8_lvt_AHMAL2
XXMn_cs_right1 vss latch_left vss latch_right sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMn_diode_right vss latch_right vss latch_right sky130_fd_pr__nfet_01v8_lvt_AHMAL2
Xsky130_fd_pr__pfet_01v8_lvt_5VNMZ8_0 out_left vdd vdd out_left vss sky130_fd_pr__pfet_01v8_lvt_5VNMZ8
XXMn_out_left vss out_left vss latch_left sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMn_out_right vss vout vss latch_right sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMp_tail tail vbias_p vdd vdd vss sky130_fd_pr__pfet_01v8_lvt_GUWLND
X0 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X1 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X2 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X3 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X4 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X5 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X6 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X7 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
C0 vbias_p out_left 0.841523f
C1 vbias_p tail 0.651669f
C2 vout vdd 1.629186f
C3 latch_right vdd 1.446106f
C4 vinp vdd 4.263518f
C5 latch_right vout 0.728353f
C6 vinn vdd 2.304739f
C7 vinp vout 0.03655f
C8 latch_left vdd 1.397101f
C9 vinn vout 0.12978f
C10 vinp latch_right 0.513108f
C11 latch_left vout 0.140137f
C12 vinn latch_right 3.535073f
C13 vinn vinp 1.25697f
C14 latch_left latch_right 5.157924f
C15 vdd out_left 2.997078f
C16 vinp latch_left 0.504304f
C17 vinn latch_left 1.33911f
C18 tail vdd 2.229149f
C19 vout out_left 0.605798f
C20 vbias_p vdd 2.119612f
C21 tail vout 0.008029f
C22 latch_right out_left 0.143102f
C23 vbias_p vout 0.144263f
C24 vinp out_left 0.225137f
C25 tail latch_right 8.894202f
C26 vinn out_left 0.081834f
C27 vbias_p latch_right 0.001093f
C28 tail vinp 2.917567f
C29 tail vinn 0.826947f
C30 vbias_p vinp 0.030109f
C31 latch_left out_left 0.73463f
C32 vbias_p vinn 0.002221f
C33 tail latch_left 8.829929f
C34 vbias_p latch_left 0.001028f
C35 tail out_left 0.006519f
C36 vinp vss 0.4258f
C37 vinn vss 0.505665f
C38 tail vss 1.097737f
C39 vbias_p vss 0.829052f
C40 vdd vss 43.54159f
C41 vout vss 3.238105f
C42 latch_right vss 4.747994f
C43 latch_left vss 5.117222f
C44 out_left vss 3.384084f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_NVJ7JE a_221_n1088# a_n163_n1088# a_n451_n1174#
+ a_n221_n1000# a_35_n1000# a_291_n1000# a_n291_n1088# a_n349_n1000# a_n35_n1088#
+ a_93_n1088# a_163_n1000# a_n93_n1000#
X0 a_163_n1000# a_93_n1088# a_35_n1000# a_n451_n1174# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X1 a_n93_n1000# a_n163_n1088# a_n221_n1000# a_n451_n1174# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X2 a_291_n1000# a_221_n1088# a_163_n1000# a_n451_n1174# sky130_fd_pr__nfet_01v8_lvt ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.35
X3 a_n221_n1000# a_n291_n1088# a_n349_n1000# a_n451_n1174# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.35
X4 a_35_n1000# a_n35_n1088# a_n93_n1000# a_n451_n1174# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
C0 a_n291_n1088# a_n349_n1000# 0.092697f
C1 a_35_n1000# a_n35_n1088# 0.092697f
C2 a_n35_n1088# a_n163_n1088# 0.104496f
C3 a_n221_n1000# a_n163_n1088# 0.092697f
C4 a_163_n1000# a_93_n1088# 0.092697f
C5 a_35_n1000# a_n93_n1000# 1.09724f
C6 a_n163_n1088# a_n93_n1000# 0.092697f
C7 a_35_n1000# a_93_n1088# 0.092697f
C8 a_n291_n1088# a_n163_n1088# 0.104496f
C9 a_35_n1000# a_163_n1000# 1.09724f
C10 a_163_n1000# a_291_n1000# 1.09724f
C11 a_221_n1088# a_93_n1088# 0.104496f
C12 a_163_n1000# a_221_n1088# 0.092697f
C13 a_n349_n1000# a_n221_n1000# 1.09724f
C14 a_n35_n1088# a_n93_n1000# 0.092697f
C15 a_n35_n1088# a_93_n1088# 0.104496f
C16 a_n221_n1000# a_n93_n1000# 1.09724f
C17 a_221_n1088# a_291_n1000# 0.092697f
C18 a_n291_n1088# a_n221_n1000# 0.092697f
C19 a_291_n1000# a_n451_n1174# 1.07603f
C20 a_163_n1000# a_n451_n1174# 0.158299f
C21 a_35_n1000# a_n451_n1174# 0.158299f
C22 a_n93_n1000# a_n451_n1174# 0.158299f
C23 a_n221_n1000# a_n451_n1174# 0.158299f
C24 a_n349_n1000# a_n451_n1174# 1.07603f
C25 a_221_n1088# a_n451_n1174# 0.308209f
C26 a_93_n1088# a_n451_n1174# 0.243769f
C27 a_n35_n1088# a_n451_n1174# 0.243694f
C28 a_n163_n1088# a_n451_n1174# 0.243769f
C29 a_n291_n1088# a_n451_n1174# 0.308209f
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_5KDBRF a_n271_n1246# a_n141_684# a_n141_n1116#
X0 a_n141_684# a_n141_n1116# a_n271_n1246# sky130_fd_pr__res_xhigh_po_1p41 l=7
C0 a_n141_684# a_n141_n1116# 0.013247f
C1 a_n141_n1116# a_n271_n1246# 0.823317f
C2 a_n141_684# a_n271_n1246# 0.823317f
.ends

.subckt timer_core V_THRESH_I DO_OUT V_DISCH_O VDD qb_sr q_sr X_SR_LATCH/X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ X_SR_LATCH/nand_0/OUT bias_3 bias_1 X_SR_LATCH/X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ v1p2 v0p6 X_SR_LATCH/nand_0/drain_mna X_COMP_P_BOTTOM/out_left bias_p V_TRIG_B_I
+ X_COMP_P_TOP/latch_left X_COMP_P_BOTTOM/latch_right out_inv3 DI_RESET_N X_COMP_P_TOP/tail
+ X_SR_LATCH/IN_R X_COMP_P_BOTTOM/tail out_inv1 VSS X_COMP_P_TOP/out_left X_COMP_P_BOTTOM/latch_left
+ X_COMP_P_TOP/latch_right X_SR_LATCH/inv_0/vout X_SR_LATCH/IN_S
XX_INV1 out_inv1 VSS VDD q_sr inv
XX_INV2[1] DO_OUT VSS VDD out_inv1 inv
XX_INV2[0] DO_OUT VSS VDD out_inv1 inv
XX_SR_LATCH X_SR_LATCH/IN_S X_SR_LATCH/IN_R DI_RESET_N q_sr VDD qb_sr X_SR_LATCH/X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ X_SR_LATCH/inv_0/vout X_SR_LATCH/nand_0/drain_mna VSS X_SR_LATCH/nand_0/OUT X_SR_LATCH/X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ sr_latch_rb
XX_COMP_P_BOTTOM v0p6 V_TRIG_B_I bias_p VDD X_COMP_P_BOTTOM/latch_left X_COMP_P_BOTTOM/tail
+ X_COMP_P_BOTTOM/out_left X_SR_LATCH/IN_S X_COMP_P_BOTTOM/latch_right VSS comp_p
XX_COMP_P_TOP V_THRESH_I v1p2 bias_p VDD X_COMP_P_TOP/latch_left X_COMP_P_TOP/tail
+ X_COMP_P_TOP/out_left X_SR_LATCH/IN_R X_COMP_P_TOP/latch_right VSS comp_p
XXMn_discharge out_inv3 out_inv3 VSS VSS VSS VSS out_inv3 V_DISCH_O out_inv3 out_inv3
+ V_DISCH_O V_DISCH_O sky130_fd_pr__nfet_01v8_lvt_NVJ7JE
XX_INV3[3] out_inv3 VSS VDD DO_OUT inv
XXR_bias_1 VSS bias_p bias_1 sky130_fd_pr__res_xhigh_po_1p41_5KDBRF
XX_INV3[2] out_inv3 VSS VDD DO_OUT inv
XXR_bias_2 VSS bias_2 bias_1 sky130_fd_pr__res_xhigh_po_1p41_5KDBRF
XX_INV3[1] out_inv3 VSS VDD DO_OUT inv
XXR_bias_3 VSS bias_2 bias_3 sky130_fd_pr__res_xhigh_po_1p41_5KDBRF
XX_INV3[0] out_inv3 VSS VDD DO_OUT inv
XXR_bias_4 VSS bias_n bias_3 sky130_fd_pr__res_xhigh_po_1p41_5KDBRF
XXR_mid VSS v0p6 v1p2 sky130_fd_pr__res_xhigh_po_1p41_5KDBRF
XXMn_bias VSS bias_n VSS bias_n sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXR_bot VSS v0p6 VSS sky130_fd_pr__res_xhigh_po_1p41_5KDBRF
XXR_top VSS VDD v1p2 sky130_fd_pr__res_xhigh_po_1p41_5KDBRF
XXMp_bias bias_p bias_p VDD VDD VSS sky130_fd_pr__pfet_01v8_lvt_GUWLND
C0 qb_sr V_DISCH_O 9.71e-19
C1 v1p2 X_SR_LATCH/IN_R 0.008984f
C2 V_DISCH_O VDD 0.009048f
C3 q_sr V_DISCH_O 7.82e-19
C4 v1p2 qb_sr 1.78e-19
C5 v1p2 VDD 1.464326f
C6 v1p2 q_sr 7.67e-21
C7 v1p2 V_THRESH_I 0.193093f
C8 v1p2 X_COMP_P_TOP/out_left 0.368388f
C9 out_inv1 V_DISCH_O 5.71e-19
C10 X_SR_LATCH/nand_0/OUT X_SR_LATCH/nand_0/drain_mna -1.91e-19
C11 X_COMP_P_TOP/tail X_COMP_P_BOTTOM/out_left 3.1e-21
C12 v1p2 out_inv1 1.53e-20
C13 X_COMP_P_BOTTOM/out_left X_COMP_P_BOTTOM/tail -0.001708f
C14 X_COMP_P_TOP/tail V_TRIG_B_I 7.62e-21
C15 bias_2 V_TRIG_B_I 0.086205f
C16 X_COMP_P_BOTTOM/out_left bias_p -0.048461f
C17 X_COMP_P_BOTTOM/tail v0p6 -0.242808f
C18 qb_sr X_SR_LATCH/nand_0/drain_mna -1.73e-19
C19 X_SR_LATCH/IN_R X_COMP_P_TOP/tail 0.002749f
C20 X_SR_LATCH/IN_R bias_2 4.01e-19
C21 bias_n V_TRIG_B_I 0.065657f
C22 X_SR_LATCH/nand_0/drain_mna VDD 0.001112f
C23 X_COMP_P_BOTTOM/tail V_TRIG_B_I -4.88e-19
C24 bias_p v0p6 -1.43e-20
C25 X_SR_LATCH/nand_0/OUT DI_RESET_N -0.016081f
C26 q_sr X_SR_LATCH/nand_0/drain_mna 2.52e-22
C27 DO_OUT X_COMP_P_BOTTOM/tail 3.93e-19
C28 bias_p V_TRIG_B_I 0.187066f
C29 bias_n X_SR_LATCH/IN_R 0.01752f
C30 DO_OUT DI_RESET_N 2.882332f
C31 DO_OUT bias_p 3.21e-19
C32 X_COMP_P_BOTTOM/out_left X_SR_LATCH/IN_S 0.574679f
C33 X_COMP_P_TOP/tail VDD 1.690042f
C34 bias_2 VDD 0.165891f
C35 X_SR_LATCH/IN_R DI_RESET_N 3.158199f
C36 X_COMP_P_TOP/tail V_THRESH_I 0.002877f
C37 X_SR_LATCH/IN_R bias_p -0.041937f
C38 V_THRESH_I bias_2 0.248813f
C39 X_SR_LATCH/IN_S v0p6 0.002374f
C40 X_SR_LATCH/nand_0/OUT X_SR_LATCH/IN_S 0.126798f
C41 bias_n VDD 0.014926f
C42 X_COMP_P_BOTTOM/out_left X_COMP_P_BOTTOM/latch_right -4.36e-19
C43 X_SR_LATCH/IN_S V_TRIG_B_I 0.009008f
C44 X_COMP_P_BOTTOM/tail VDD 2.207734f
C45 bias_n V_THRESH_I 0.252991f
C46 qb_sr DI_RESET_N -0.007459f
C47 DO_OUT X_SR_LATCH/IN_S 0.110481f
C48 DI_RESET_N VDD 0.787561f
C49 X_COMP_P_BOTTOM/latch_right v0p6 -3.54e-19
C50 bias_p VDD 4.9051f
C51 X_COMP_P_BOTTOM/tail X_COMP_P_TOP/out_left 3.1e-21
C52 q_sr DI_RESET_N -8.7e-19
C53 X_SR_LATCH/IN_R X_SR_LATCH/IN_S 0.163728f
C54 V_THRESH_I bias_p 0.069459f
C55 bias_p X_COMP_P_TOP/out_left 0.003913f
C56 X_SR_LATCH/inv_0/vout DI_RESET_N 0.003006f
C57 DO_OUT X_COMP_P_BOTTOM/latch_right 4.16e-19
C58 X_SR_LATCH/IN_S out_inv3 0.177402f
C59 qb_sr X_SR_LATCH/IN_S 0.138415f
C60 X_COMP_P_BOTTOM/out_left X_COMP_P_BOTTOM/latch_left -9.54e-19
C61 X_SR_LATCH/IN_S VDD 0.6047f
C62 q_sr X_SR_LATCH/IN_S 0.03636f
C63 DO_OUT bias_1 4.12e-19
C64 X_COMP_P_BOTTOM/latch_right out_inv3 0.003058f
C65 X_SR_LATCH/IN_S X_COMP_P_TOP/out_left 0.016125f
C66 X_SR_LATCH/inv_0/vout X_SR_LATCH/IN_S 0.004418f
C67 X_SR_LATCH/IN_R bias_1 0.005393f
C68 X_COMP_P_BOTTOM/latch_right VDD 0.248896f
C69 v1p2 X_COMP_P_TOP/tail 6.78e-20
C70 v1p2 bias_2 2.52e-19
C71 DO_OUT X_COMP_P_BOTTOM/latch_left 2.39e-19
C72 out_inv1 X_SR_LATCH/IN_S 0.046883f
C73 bias_1 VDD 0.364699f
C74 X_COMP_P_BOTTOM/latch_left out_inv3 0.029394f
C75 v1p2 DI_RESET_N 5.91e-19
C76 v1p2 bias_p 0.358806f
C77 X_COMP_P_BOTTOM/latch_left VDD 0.44241f
C78 V_DISCH_O X_SR_LATCH/IN_S 0.25997f
C79 v1p2 X_SR_LATCH/IN_S 1.61e-19
C80 DI_RESET_N X_SR_LATCH/nand_0/drain_mna 4.5e-21
C81 V_DISCH_O X_COMP_P_BOTTOM/latch_left 8.96e-20
C82 bias_n bias_2 0.069293f
C83 bias_p bias_2 0.069263f
C84 X_SR_LATCH/nand_0/drain_mna X_SR_LATCH/IN_S 0.005048f
C85 bias_p X_COMP_P_BOTTOM/tail -0.001021f
C86 DI_RESET_N bias_p 3.36e-19
C87 X_SR_LATCH/IN_S X_COMP_P_BOTTOM/tail 0.002753f
C88 DO_OUT bias_3 4.12e-19
C89 DI_RESET_N X_SR_LATCH/IN_S 0.065921f
C90 X_SR_LATCH/IN_S bias_p -0.049709f
C91 X_SR_LATCH/IN_R bias_3 0.01147f
C92 X_COMP_P_BOTTOM/latch_right X_COMP_P_BOTTOM/tail -0.001124f
C93 bias_1 bias_2 6.55e-19
C94 X_COMP_P_BOTTOM/latch_right bias_p -3.02e-19
C95 X_COMP_P_TOP/latch_left V_TRIG_B_I 2.85e-19
C96 bias_3 VDD 0.028714f
C97 DI_RESET_N bias_1 6e-19
C98 X_SR_LATCH/IN_R X_COMP_P_TOP/latch_left 0.12645f
C99 bias_1 bias_p 0.043358f
C100 X_COMP_P_BOTTOM/latch_right X_SR_LATCH/IN_S 0.168326f
C101 X_COMP_P_BOTTOM/latch_left X_COMP_P_BOTTOM/tail -0.001942f
C102 X_COMP_P_BOTTOM/latch_left bias_p -4.71e-19
C103 X_COMP_P_TOP/latch_left VDD 0.419421f
C104 X_COMP_P_TOP/latch_left V_THRESH_I 0.02646f
C105 X_COMP_P_BOTTOM/latch_left X_SR_LATCH/IN_S 0.122408f
C106 X_COMP_P_TOP/latch_right V_TRIG_B_I 4.9e-21
C107 X_COMP_P_BOTTOM/out_left v0p6 0.008241f
C108 v1p2 X_COMP_P_TOP/latch_left 3.97e-20
C109 X_COMP_P_BOTTOM/out_left V_TRIG_B_I 0.300686f
C110 X_SR_LATCH/IN_R X_COMP_P_TOP/latch_right 0.128018f
C111 DO_OUT X_COMP_P_BOTTOM/out_left 0.13262f
C112 V_TRIG_B_I v0p6 0.112639f
C113 X_SR_LATCH/IN_R X_COMP_P_BOTTOM/out_left 0.016095f
C114 X_SR_LATCH/X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# out_inv3 1.51e-20
C115 DO_OUT v0p6 0.431659f
C116 DO_OUT X_SR_LATCH/nand_0/OUT 7.62e-19
C117 X_COMP_P_TOP/latch_right VDD 0.212823f
C118 X_SR_LATCH/X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# VDD 0.011923f
C119 DO_OUT V_TRIG_B_I 0.347624f
C120 X_COMP_P_BOTTOM/out_left out_inv3 0.013941f
C121 X_COMP_P_TOP/latch_right V_THRESH_I 0.002476f
C122 q_sr X_SR_LATCH/X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 0.001244f
C123 X_SR_LATCH/X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# VDD 0.011952f
C124 X_SR_LATCH/IN_R V_TRIG_B_I 0.084879f
C125 X_COMP_P_BOTTOM/out_left VDD 1.202144f
C126 out_inv3 v0p6 0.002838f
C127 q_sr X_SR_LATCH/X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# 0.003779f
C128 X_SR_LATCH/IN_R DO_OUT 0.060174f
C129 X_COMP_P_BOTTOM/out_left V_THRESH_I 1e-20
C130 X_SR_LATCH/nand_0/OUT out_inv3 1.61e-19
C131 bias_3 bias_2 6.55e-19
C132 X_COMP_P_BOTTOM/out_left X_COMP_P_TOP/out_left 0.016634f
C133 X_SR_LATCH/nand_0/OUT qb_sr -1.49e-19
C134 out_inv3 V_TRIG_B_I 0.217319f
C135 VDD v0p6 1.67662f
C136 X_SR_LATCH/nand_0/OUT VDD 0.06012f
C137 DO_OUT out_inv3 0.667717f
C138 X_COMP_P_TOP/out_left v0p6 6.4e-22
C139 VDD V_TRIG_B_I 1.079768f
C140 DO_OUT qb_sr 8.53e-19
C141 q_sr X_SR_LATCH/nand_0/OUT 0.024468f
C142 bias_n bias_3 6.55e-19
C143 DO_OUT VDD 1.810194f
C144 V_THRESH_I V_TRIG_B_I 0.565173f
C145 X_SR_LATCH/nand_0/OUT X_SR_LATCH/inv_0/vout -1.88e-19
C146 X_COMP_P_TOP/out_left V_TRIG_B_I 0.144366f
C147 q_sr DO_OUT 7.86e-20
C148 out_inv1 X_COMP_P_BOTTOM/out_left 1.75e-19
C149 DI_RESET_N bias_3 6e-19
C150 bias_3 bias_p 6.09e-20
C151 X_SR_LATCH/IN_R VDD 1.592842f
C152 DO_OUT X_SR_LATCH/inv_0/vout 4.72e-20
C153 q_sr X_SR_LATCH/IN_R 0.001378f
C154 X_SR_LATCH/IN_R V_THRESH_I 0.063976f
C155 qb_sr out_inv3 6.26e-19
C156 X_SR_LATCH/IN_R X_COMP_P_TOP/out_left 0.396136f
C157 X_SR_LATCH/IN_R X_SR_LATCH/inv_0/vout 0.005005f
C158 VDD out_inv3 0.643841f
C159 out_inv1 X_SR_LATCH/nand_0/OUT 0.001405f
C160 qb_sr VDD 0.040093f
C161 q_sr out_inv3 2.38e-20
C162 q_sr qb_sr 0.004823f
C163 bias_n X_COMP_P_TOP/latch_left 0.001099f
C164 out_inv1 DO_OUT 0.35078f
C165 q_sr VDD 0.275245f
C166 V_THRESH_I VDD 0.935463f
C167 X_SR_LATCH/inv_0/vout qb_sr -8.15e-20
C168 v1p2 X_COMP_P_TOP/latch_right 2.09e-20
C169 X_COMP_P_TOP/out_left VDD 1.184775f
C170 out_inv1 X_SR_LATCH/IN_R 3.82e-22
C171 X_SR_LATCH/inv_0/vout VDD 0.025978f
C172 V_THRESH_I X_COMP_P_TOP/out_left 0.017536f
C173 q_sr X_SR_LATCH/inv_0/vout 2.81e-19
C174 X_SR_LATCH/nand_0/OUT V_DISCH_O 0.00105f
C175 v1p2 X_COMP_P_BOTTOM/out_left 0.008724f
C176 out_inv1 qb_sr 0.002285f
C177 DO_OUT V_DISCH_O 8.56e-19
C178 v1p2 v0p6 0.158301f
C179 out_inv1 VDD 0.313959f
C180 v1p2 X_SR_LATCH/nand_0/OUT 1.51e-19
C181 out_inv1 q_sr 0.160379f
C182 bias_3 bias_1 0.06887f
C183 v1p2 V_TRIG_B_I 1.116621f
C184 out_inv1 X_SR_LATCH/inv_0/vout 1.05e-20
C185 v1p2 DO_OUT 0.150366f
C186 V_DISCH_O out_inv3 0.326617f
C187 v1p2 VSS 3.146392f
C188 bias_n VSS 2.376644f
C189 bias_3 VSS 1.654247f
C190 bias_2 VSS 1.434531f
C191 bias_1 VSS 1.576978f
C192 VDD VSS 99.65678f
C193 DO_OUT VSS 2.622944f
C194 V_DISCH_O VSS 5.743176f
C195 out_inv3 VSS 3.448332f
C196 V_THRESH_I VSS 1.49496f
C197 X_COMP_P_TOP/tail VSS 1.14054f
C198 X_COMP_P_TOP/latch_right VSS 4.224772f
C199 X_COMP_P_TOP/latch_left VSS 3.910736f
C200 X_COMP_P_TOP/out_left VSS 2.068422f
C201 v0p6 VSS 2.245097f
C202 V_TRIG_B_I VSS 1.423111f
C203 X_COMP_P_BOTTOM/tail VSS 1.140396f
C204 bias_p VSS 2.867893f
C205 X_SR_LATCH/IN_S VSS 8.636353f
C206 X_COMP_P_BOTTOM/latch_right VSS 4.31988f
C207 X_COMP_P_BOTTOM/latch_left VSS 3.964322f
C208 X_COMP_P_BOTTOM/out_left VSS 2.072656f
C209 X_SR_LATCH/nand_0/drain_mna VSS 0.108699f
C210 X_SR_LATCH/nand_0/OUT VSS 0.531925f
C211 DI_RESET_N VSS 1.742971f
C212 qb_sr VSS 0.560008f
C213 X_SR_LATCH/X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# VSS 0.020511f
C214 X_SR_LATCH/X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# VSS 0.020511f
C215 X_SR_LATCH/inv_0/vout VSS 0.394084f
C216 X_SR_LATCH/IN_R VSS 11.2019f
C217 out_inv1 VSS 0.672412f
C218 q_sr VSS 0.826371f
.ends

.subckt tt_um_vaf_555_timer clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VPWR VGND
XX_TIMER ua[0] uo_out[0] ua[2] VPWR X_TIMER/qb_sr X_TIMER/q_sr X_TIMER/X_SR_LATCH/X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ X_TIMER/X_SR_LATCH/nand_0/OUT X_TIMER/bias_3 X_TIMER/bias_1 X_TIMER/X_SR_LATCH/X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164#
+ X_TIMER/v1p2 X_TIMER/v0p6 X_TIMER/X_SR_LATCH/nand_0/drain_mna X_TIMER/X_COMP_P_BOTTOM/out_left
+ X_TIMER/bias_p ua[1] X_TIMER/X_COMP_P_TOP/latch_left X_TIMER/X_COMP_P_BOTTOM/latch_right
+ X_TIMER/out_inv3 ui_in[0] X_TIMER/X_COMP_P_TOP/tail X_TIMER/X_SR_LATCH/IN_R X_TIMER/X_COMP_P_BOTTOM/tail
+ X_TIMER/out_inv1 VGND X_TIMER/X_COMP_P_TOP/out_left X_TIMER/X_COMP_P_BOTTOM/latch_left
+ X_TIMER/X_COMP_P_TOP/latch_right X_TIMER/X_SR_LATCH/inv_0/vout X_TIMER/X_SR_LATCH/IN_S
+ timer_core
C0 X_TIMER/qb_sr ua[2] 1.66e-20
C1 ua[1] X_TIMER/v0p6 0.009908f
C2 uo_out[0] uio_oe[1] 0.013858f
C3 ua[3] ua[2] 0.0564f
C4 uio_out[4] uio_out[3] 0.023797f
C5 ua[4] ua[2] 0.0564f
C6 ua[5] ua[2] 0.0564f
C7 uio_in[6] uio_in[5] 0.023797f
C8 uo_out[0] uo_out[7] 0.013858f
C9 X_TIMER/X_COMP_P_BOTTOM/out_left ua[2] 0.005338f
C10 X_TIMER/out_inv1 VPWR 1.26e-20
C11 uio_out[0] uo_out[0] 0.013858f
C12 uio_in[4] uio_in[5] 0.023797f
C13 uo_out[0] uio_oe[5] 0.013858f
C14 uio_oe[0] uio_out[7] 0.023797f
C15 uo_out[0] uo_out[6] 0.013858f
C16 uio_oe[1] uio_oe[2] 0.023797f
C17 uio_in[4] uio_in[3] 0.023797f
C18 X_TIMER/X_SR_LATCH/X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# VPWR 0.001066f
C19 uio_in[5] ui_in[0] 0.010273f
C20 uio_in[6] ui_in[0] 0.010273f
C21 ui_in[0] VPWR 0.246688f
C22 uio_in[3] ui_in[0] 0.010273f
C23 uio_oe[3] uio_oe[4] 0.023797f
C24 X_TIMER/X_SR_LATCH/IN_R ua[0] 0.031154f
C25 uio_in[4] ui_in[0] 0.010273f
C26 ui_in[3] ui_in[2] 0.023797f
C27 uo_out[2] uo_out[1] 0.023797f
C28 ui_in[6] ui_in[7] 0.023797f
C29 X_TIMER/v1p2 ua[1] 0.007859f
C30 X_TIMER/X_COMP_P_TOP/latch_left ua[0] 0.002454f
C31 uio_in[6] uio_in[7] 0.023797f
C32 uo_out[0] uo_out[1] 0.037655f
C33 X_TIMER/X_COMP_P_BOTTOM/tail ua[1] 0.01003f
C34 clk ena 0.023797f
C35 ua[2] VPWR 0.025379f
C36 X_TIMER/X_COMP_P_TOP/out_left ua[0] 0.002039f
C37 uio_oe[0] uo_out[0] 0.013858f
C38 uio_out[0] uio_out[1] 0.023797f
C39 ua[2] X_TIMER/X_COMP_P_BOTTOM/latch_left 0.011668f
C40 ui_in[0] uio_in[7] 0.010273f
C41 uio_out[7] uio_out[6] 0.023797f
C42 ua[1] ua[0] 10.177747f
C43 uo_out[0] VPWR 5.339137f
C44 X_TIMER/X_COMP_P_BOTTOM/out_left ua[1] 0.006774f
C45 uo_out[0] uio_oe[4] 0.013858f
C46 uo_out[5] uo_out[0] 0.013858f
C47 uio_oe[6] uo_out[0] 0.013858f
C48 uo_out[0] uio_oe[3] 0.013858f
C49 uio_out[7] uo_out[0] 0.013858f
C50 X_TIMER/X_SR_LATCH/IN_R VPWR 0.1463f
C51 ui_in[0] uo_out[0] 16.853556f
C52 X_TIMER/X_SR_LATCH/IN_S VPWR 0.020214f
C53 ui_in[0] ui_in[1] 0.034283f
C54 ui_in[0] ui_in[2] 0.010273f
C55 ui_in[6] ui_in[5] 0.023797f
C56 uo_out[0] uio_in[7] 0.023797f
C57 X_TIMER/X_SR_LATCH/nand_0/drain_mna VPWR 0.001225f
C58 ui_in[0] X_TIMER/X_SR_LATCH/IN_R 0.045844f
C59 uio_out[6] uo_out[0] 0.013858f
C60 X_TIMER/X_SR_LATCH/X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# VPWR 0.001585f
C61 uio_out[0] uo_out[7] 0.023797f
C62 uio_oe[3] uio_oe[2] 0.023797f
C63 X_TIMER/bias_3 VPWR 0.02155f
C64 ua[1] VPWR 0.17723f
C65 uio_in[3] uio_in[2] 0.023797f
C66 X_TIMER/q_sr VPWR 0.006835f
C67 ui_in[0] rst_n 0.02398f
C68 ua[1] X_TIMER/X_COMP_P_TOP/tail 0.010049f
C69 uo_out[7] uo_out[6] 0.023797f
C70 uio_oe[6] uio_oe[7] 0.023797f
C71 uo_out[0] uo_out[2] 0.013858f
C72 ui_in[0] ui_in[7] 0.010273f
C73 X_TIMER/out_inv3 VPWR 0.004294f
C74 uio_out[6] uio_out[5] 0.023797f
C75 ui_in[5] ui_in[4] 0.023797f
C76 ui_in[0] uio_in[0] 0.010273f
C77 ua[1] X_TIMER/X_COMP_P_BOTTOM/latch_left 0.015471f
C78 ui_in[0] uio_in[1] 0.010273f
C79 uo_out[5] uo_out[4] 0.023797f
C80 ua[2] X_TIMER/X_SR_LATCH/IN_S 0.014944f
C81 ui_in[0] uio_in[2] 0.010273f
C82 ua[1] X_TIMER/X_COMP_P_TOP/latch_right 0.090134f
C83 ua[2] X_TIMER/X_COMP_P_BOTTOM/latch_right 0.011181f
C84 uo_out[0] X_TIMER/X_SR_LATCH/IN_R 1.12e-19
C85 X_TIMER/X_SR_LATCH/nand_0/OUT VPWR 0.011264f
C86 uo_out[0] uio_out[5] 0.013858f
C87 uio_oe[0] uio_oe[1] 0.023797f
C88 ui_in[2] ui_in[1] 0.023797f
C89 uio_out[2] uo_out[0] 0.013858f
C90 uo_out[0] uio_oe[2] 0.013858f
C91 uo_out[2] uo_out[3] 0.023797f
C92 ua[1] ua[2] 4.93575f
C93 ui_in[4] ui_in[3] 0.023797f
C94 ua[2] X_TIMER/q_sr 1.17e-20
C95 uo_out[0] uo_out[3] 0.013858f
C96 X_TIMER/bias_1 VPWR 0.022502f
C97 X_TIMER/v1p2 VPWR 0.044876f
C98 X_TIMER/out_inv3 ua[2] 0.012327f
C99 uio_out[4] uo_out[0] 0.013858f
C100 X_TIMER/bias_p VPWR 0.033435f
C101 uo_out[0] uo_out[4] 0.013858f
C102 uo_out[0] uio_out[1] 0.013858f
C103 X_TIMER/X_SR_LATCH/nand_0/OUT ua[2] 1.66e-20
C104 X_TIMER/qb_sr VPWR 0.005282f
C105 uo_out[0] uio_out[3] 0.013858f
C106 ua[7] VPWR 0.010285f
C107 ui_in[5] ui_in[0] 0.010273f
C108 X_TIMER/X_SR_LATCH/inv_0/vout VPWR 0.01271f
C109 uio_out[4] uio_out[5] 0.023797f
C110 rst_n clk 0.023797f
C111 ui_in[6] ui_in[0] 0.010273f
C112 uio_oe[5] uio_oe[4] 0.023797f
C113 X_TIMER/X_SR_LATCH/IN_R ua[1] 0.051759f
C114 X_TIMER/X_COMP_P_TOP/latch_left ua[1] 0.070843f
C115 ua[1] X_TIMER/X_SR_LATCH/IN_S 0.006697f
C116 uio_oe[6] uio_oe[5] 0.023797f
C117 uo_out[5] uo_out[6] 0.023797f
C118 uio_out[2] uio_out[1] 0.023797f
C119 ua[1] X_TIMER/X_COMP_P_BOTTOM/latch_right 0.040903f
C120 uio_in[0] ui_in[7] 0.023797f
C121 uo_out[3] uo_out[4] 0.023797f
C122 uio_out[2] uio_out[3] 0.023797f
C123 X_TIMER/X_COMP_P_TOP/latch_right ua[0] 2.47e-19
C124 X_TIMER/X_COMP_P_TOP/out_left ua[1] 0.016671f
C125 uio_in[0] uio_in[1] 0.023797f
C126 ui_in[0] ui_in[3] 0.010273f
C127 uio_in[2] uio_in[1] 0.023797f
C128 ui_in[0] ui_in[4] 0.010273f
C129 ua[2] ua[6] 0.0564f
C130 ua[3] VGND 0.101433f
C131 ua[4] VGND 0.101433f
C132 ua[5] VGND 0.101909f
C133 ua[6] VGND 0.102993f
C134 ua[7] VGND 0.112606f
C135 ena VGND 0.073297f
C136 clk VGND 0.0487f
C137 rst_n VGND 0.04861f
C138 ui_in[1] VGND 0.040051f
C139 ui_in[2] VGND 0.040155f
C140 ui_in[3] VGND 0.040155f
C141 ui_in[4] VGND 0.040155f
C142 ui_in[5] VGND 0.040155f
C143 ui_in[6] VGND 0.040155f
C144 ui_in[7] VGND 0.040155f
C145 uio_in[0] VGND 0.040155f
C146 uio_in[1] VGND 0.040155f
C147 uio_in[2] VGND 0.040155f
C148 uio_in[3] VGND 0.040155f
C149 uio_in[4] VGND 0.040155f
C150 uio_in[5] VGND 0.040155f
C151 uio_in[6] VGND 0.040155f
C152 uio_in[7] VGND 0.040155f
C153 uo_out[1] VGND 0.03939f
C154 uo_out[2] VGND 0.03939f
C155 uo_out[3] VGND 0.03939f
C156 uo_out[4] VGND 0.03939f
C157 uo_out[5] VGND 0.03939f
C158 uo_out[6] VGND 0.03939f
C159 uo_out[7] VGND 0.03939f
C160 uio_out[0] VGND 0.03939f
C161 uio_out[1] VGND 0.03939f
C162 uio_out[2] VGND 0.03939f
C163 uio_out[3] VGND 0.03939f
C164 uio_out[4] VGND 0.03939f
C165 uio_out[5] VGND 0.03939f
C166 uio_out[6] VGND 0.03939f
C167 uio_out[7] VGND 0.03939f
C168 uio_oe[0] VGND 0.03939f
C169 uio_oe[1] VGND 0.03939f
C170 uio_oe[2] VGND 0.03939f
C171 uio_oe[3] VGND 0.03939f
C172 uio_oe[4] VGND 0.03939f
C173 uio_oe[5] VGND 0.03939f
C174 uio_oe[6] VGND 0.03939f
C175 uio_oe[7] VGND 0.073297f
C176 X_TIMER/v1p2 VGND 2.527758f
C177 X_TIMER/bias_n VGND 1.931379f
C178 X_TIMER/bias_3 VGND 1.580737f
C179 X_TIMER/bias_2 VGND 1.393845f
C180 X_TIMER/bias_1 VGND 1.521669f
C181 VPWR VGND 0.108412p
C182 uo_out[0] VGND 9.090312f
C183 ua[2] VGND 7.393198f
C184 X_TIMER/out_inv3 VGND 2.186164f
C185 ua[0] VGND 16.42065f
C186 X_TIMER/X_COMP_P_TOP/tail VGND 1.097679f
C187 X_TIMER/X_COMP_P_TOP/latch_right VGND 3.519466f
C188 X_TIMER/X_COMP_P_TOP/latch_left VGND 3.688133f
C189 X_TIMER/X_COMP_P_TOP/out_left VGND 2.066467f
C190 X_TIMER/v0p6 VGND 2.033237f
C191 ua[1] VGND 11.711487f
C192 X_TIMER/X_COMP_P_BOTTOM/tail VGND 1.097675f
C193 X_TIMER/bias_p VGND 2.785426f
C194 X_TIMER/X_SR_LATCH/IN_S VGND 2.669827f
C195 X_TIMER/X_COMP_P_BOTTOM/latch_right VGND 3.519416f
C196 X_TIMER/X_COMP_P_BOTTOM/latch_left VGND 3.688127f
C197 X_TIMER/X_COMP_P_BOTTOM/out_left VGND 2.066463f
C198 X_TIMER/X_SR_LATCH/nand_0/drain_mna VGND 0.108169f
C199 X_TIMER/X_SR_LATCH/nand_0/OUT VGND 0.524253f
C200 ui_in[0] VGND 16.823254f
C201 X_TIMER/qb_sr VGND 0.53504f
C202 X_TIMER/X_SR_LATCH/X_NOR_BOTTOM/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# VGND 0.020446f
C203 X_TIMER/X_SR_LATCH/X_NOR_TOP/sky130_fd_pr__pfet_01v8_7P3MHC_1/a_14_n164# VGND 0.020446f
C204 X_TIMER/X_SR_LATCH/inv_0/vout VGND 0.337759f
C205 X_TIMER/X_SR_LATCH/IN_R VGND 3.018241f
C206 X_TIMER/out_inv1 VGND 0.5524f
C207 X_TIMER/q_sr VGND 0.736573f
.ends

