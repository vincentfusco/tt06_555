magic
tech sky130A
magscale 1 2
timestamp 1711739992
<< nwell >>
rect 23452 19652 23920 20064
rect 20680 18281 23158 18315
<< pwell >>
rect 20680 17271 23166 17305
<< psubdiff >>
rect 20680 17271 23166 17305
<< nsubdiff >>
rect 24102 19798 28001 19916
rect 20680 18281 23158 18315
<< locali >>
rect 23452 19916 23920 20064
rect 23402 19798 28613 19916
rect 23452 19652 23920 19798
<< viali >>
rect 20810 20140 22984 20174
<< metal1 >>
rect 20631 23478 20641 23878
rect 28516 23478 28587 23878
rect 25275 20548 25285 20604
rect 25661 20548 25671 20604
rect 26475 20548 26485 20604
rect 26861 20548 26871 20604
rect 20800 20180 20810 20184
rect 20798 20134 20810 20180
rect 22984 20180 22994 20184
rect 20800 20132 20810 20134
rect 22984 20134 22996 20180
rect 22984 20132 22994 20134
rect 23452 19916 23920 20064
rect 23402 19798 23522 19916
rect 28577 19798 28613 19916
rect 23452 19652 23920 19798
rect 25275 19110 25285 19166
rect 25661 19110 25671 19166
rect 26475 19110 26485 19166
rect 26861 19110 26871 19166
rect 24432 18538 24442 18590
rect 25395 18538 25405 18590
rect 20646 18281 20656 18333
rect 23181 18281 23191 18333
rect 20680 17271 23166 17305
rect 20810 16448 20856 17030
rect 22920 16448 22966 17030
rect 20678 16276 28610 16338
rect 20678 16236 28614 16276
rect 20667 15836 20677 16236
rect 28613 15836 28623 16236
<< via1 >>
rect 20641 23478 28516 23878
rect 25285 20548 25661 20604
rect 26485 20548 26861 20604
rect 20810 20174 22984 20184
rect 20810 20140 22984 20174
rect 20810 20132 22984 20140
rect 23522 19798 28577 19916
rect 25285 19110 25661 19166
rect 26485 19110 26861 19166
rect 24442 18538 25395 18590
rect 20656 18281 23181 18333
rect 20677 15836 28613 16236
<< metal2 >>
rect 20641 23878 28577 23888
rect 28516 23478 28578 23878
rect 20641 23468 28577 23478
rect 25285 20604 25661 20614
rect 25285 20538 25661 20548
rect 26485 20604 26861 20614
rect 26485 20538 26861 20548
rect 20810 20184 22984 20194
rect 20810 20068 22984 20132
rect 28000 20068 28613 20069
rect 20428 20058 28613 20068
rect 20428 19916 24103 20058
rect 27308 19916 28613 20058
rect 20428 19798 23522 19916
rect 28577 19798 28613 19916
rect 20428 19658 24103 19798
rect 27308 19658 28613 19798
rect 20428 19648 28613 19658
rect 25285 19166 25661 19176
rect 25285 19100 25661 19110
rect 26485 19166 26861 19176
rect 26485 19100 26861 19110
rect 24442 18594 25395 18604
rect 24442 18528 25395 18538
rect 20656 18337 23181 18347
rect 20656 18271 23181 18281
rect 20677 16236 28613 16246
rect 20677 15826 28613 15836
<< via2 >>
rect 20641 23478 28166 23878
rect 25285 20548 25661 20604
rect 26485 20548 26861 20604
rect 24103 19916 27308 20058
rect 24103 19798 27308 19916
rect 24103 19658 27308 19798
rect 25285 19110 25661 19166
rect 26485 19110 26861 19166
rect 24442 18590 25395 18594
rect 24442 18538 25395 18590
rect 20656 18333 23181 18337
rect 20656 18281 23181 18333
rect 20677 15836 28166 16236
<< metal3 >>
rect 20631 23878 28613 23883
rect 20631 23874 20641 23878
rect 20428 23478 20641 23874
rect 28166 23478 28613 23878
rect 20428 23474 28613 23478
rect 20631 23473 28613 23474
rect 20428 21123 26861 21523
rect 25285 20609 25661 21123
rect 26485 20609 26861 21123
rect 25275 20604 25671 20609
rect 25275 20548 25285 20604
rect 25661 20548 25671 20604
rect 25275 20543 25671 20548
rect 26475 20604 26871 20609
rect 26475 20548 26485 20604
rect 26861 20548 26871 20604
rect 26475 20543 26871 20548
rect 20428 20063 24103 20068
rect 25285 20063 25661 20543
rect 26485 20063 26861 20543
rect 27308 20063 27568 20068
rect 20428 20058 27568 20063
rect 20428 19658 24103 20058
rect 27308 19658 27568 20058
rect 20428 19653 27568 19658
rect 20428 19648 24103 19653
rect 25285 19171 25661 19653
rect 26485 19171 26861 19653
rect 27308 19648 27568 19653
rect 25275 19166 25671 19171
rect 25275 19110 25285 19166
rect 25661 19110 25671 19166
rect 25275 19105 25671 19110
rect 26475 19166 26871 19171
rect 26475 19110 26485 19166
rect 26861 19110 26871 19166
rect 26475 19105 26871 19110
rect 25285 18599 25661 19105
rect 24432 18594 25661 18599
rect 24432 18592 24442 18594
rect 20428 18538 24442 18592
rect 25395 18592 25661 18594
rect 26485 18630 26861 19105
rect 26485 18592 26860 18630
rect 25395 18538 26860 18592
rect 20428 18337 26860 18538
rect 20428 18281 20656 18337
rect 23181 18281 26860 18337
rect 20428 18192 26860 18281
rect 28213 16241 28613 23473
rect 20667 16236 28613 16241
rect 20667 16231 20677 16236
rect 20428 15836 20677 16231
rect 28166 15894 28613 16236
rect 28166 15836 28623 15894
rect 20428 15831 28623 15836
use comp_p  X_COMP_P_BOTTOM
timestamp 1711732688
transform 1 0 26492 0 1 14702
box -3002 1462 2120 5166
use comp_p  X_COMP_P_TOP
timestamp 1711732688
transform 1 0 26493 0 -1 25012
box -3002 1462 2120 5166
use inv  X_INV1
timestamp 1711732688
transform 1 0 20381 0 1 16477
box 978 788 1260 1874
use inv  X_INV2[0]
timestamp 1711732688
transform 1 0 20906 0 1 16477
box 978 788 1260 1874
use inv  X_INV2[1]
timestamp 1711732688
transform 1 0 20643 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[0]
timestamp 1711732688
transform 1 0 21958 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[1]
timestamp 1711732688
transform 1 0 21695 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[2]
timestamp 1711732688
transform 1 0 21432 0 1 16477
box 978 788 1260 1874
use inv  X_INV3[3]
timestamp 1711732688
transform 1 0 21169 0 1 16477
box 978 788 1260 1874
use sr_latch  X_SR_LATCH
timestamp 1711732688
transform -1 0 15343 0 1 16911
box -6020 354 -5267 1440
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_bias
timestamp 1711732688
transform 0 1 21906 -1 0 23184
box -296 -734 296 766
use sky130_fd_pr__nfet_01v8_lvt_NVJ7JE  XMn_discharge
timestamp 1711736161
transform 0 1 21888 -1 0 16739
box -487 -1210 487 1210
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_bias
timestamp 1711732688
transform 0 1 21897 -1 0 20400
box -296 -1219 296 1219
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_1
timestamp 1711732688
transform 0 1 21914 1 0 21055
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_2
timestamp 1711732688
transform 0 1 21914 1 0 21563
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_3
timestamp 1711732688
transform 0 1 21914 1 0 22071
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_4
timestamp 1711732688
transform 0 1 21914 1 0 22579
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bot
timestamp 1711732688
transform 0 1 21914 -1 0 18731
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_mid
timestamp 1711732688
transform 0 1 21914 -1 0 19239
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_top
timestamp 1711732688
transform 0 1 21914 -1 0 19747
box -307 -1282 307 1282
<< end >>
