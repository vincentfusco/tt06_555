magic
tech sky130A
magscale 1 2
timestamp 1711683265
<< error_p >>
rect 4726 14974 4772 14986
rect 5254 14974 5300 14986
rect 4726 14940 4732 14974
rect 5254 14940 5260 14974
rect 4726 14928 4772 14940
rect 5254 14928 5300 14940
rect 4726 14658 4772 14670
rect 5254 14658 5300 14670
rect 4726 14624 4732 14658
rect 5254 14624 5260 14658
rect 4726 14612 4772 14624
rect 5254 14612 5300 14624
rect 4826 14200 4872 14212
rect 5136 14200 5182 14212
rect 4826 14166 4832 14200
rect 5136 14166 5142 14200
rect 4826 14154 4872 14166
rect 5136 14154 5182 14166
rect 4826 13884 4872 13896
rect 5136 13884 5182 13896
rect 4826 13850 4832 13884
rect 5136 13850 5142 13884
rect 4826 13838 4872 13850
rect 5136 13838 5182 13850
<< error_s >>
rect 24103 19882 28001 19886
rect 30565 18344 30569 18797
rect 30593 18344 30597 18797
rect 30565 18139 30569 18168
rect 30593 18167 30597 18168
rect 30922 18167 30943 18973
rect 30950 18567 31197 19205
rect 30950 18139 30971 18567
rect 31351 18167 31372 18973
rect 31379 18567 31626 19205
rect 31379 18139 31400 18567
rect 31780 18167 31801 18973
rect 31808 18567 32055 19205
rect 31808 18139 31829 18567
rect 32209 18167 32230 18973
rect 32237 18567 32484 19205
rect 32237 18139 32258 18567
rect 32638 18167 32659 18973
rect 32666 18567 32913 19205
rect 32666 18139 32687 18567
<< error_ps >>
rect 11400 19292 11446 19304
rect 11928 19292 11974 19304
rect 11400 19258 11406 19292
rect 11928 19258 11934 19292
rect 11400 19246 11446 19258
rect 11928 19246 11974 19258
rect 11400 18976 11446 18988
rect 11928 18976 11974 18988
rect 11400 18942 11406 18976
rect 11928 18942 11934 18976
rect 11400 18930 11446 18942
rect 11928 18930 11974 18942
rect 11500 18518 11546 18530
rect 11810 18518 11856 18530
rect 11500 18484 11506 18518
rect 11810 18484 11816 18518
rect 11500 18472 11546 18484
rect 11810 18472 11856 18484
rect 11500 18202 11546 18214
rect 11810 18202 11856 18214
rect 11500 18168 11506 18202
rect 11810 18168 11816 18202
rect 11500 18156 11546 18168
rect 11810 18156 11856 18168
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use comp_p  comp_p_0
timestamp 1711658383
transform 1 0 26493 0 -1 25012
box -3002 1462 2120 5166
use comp_p  X_COMP_P1
timestamp 1711658383
transform 1 0 26492 0 1 14702
box -3002 1462 2120 5166
use inv  X_INV1
timestamp 1711045747
transform 1 0 30265 0 1 17385
box -60 547 369 1820
use inv  X_INV2[0]
timestamp 1711045747
transform 1 0 31010 0 1 17385
box -60 547 369 1820
use inv  X_INV2[1]
timestamp 1711045747
transform 1 0 30581 0 1 17385
box -60 547 369 1820
use inv  X_INV3[0]
timestamp 1711045747
transform 1 0 32726 0 1 17385
box -60 547 369 1820
use inv  X_INV3[1]
timestamp 1711045747
transform 1 0 32297 0 1 17385
box -60 547 369 1820
use inv  X_INV3[2]
timestamp 1711045747
transform 1 0 31868 0 1 17385
box -60 547 369 1820
use inv  X_INV3[3]
timestamp 1711045747
transform 1 0 31439 0 1 17385
box -60 547 369 1820
use sr_latch  X_SR_LATCH
timestamp 1711045747
transform 1 0 8745 0 1 14056
box -4457 -2000 3703 5706
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XMn_bias
timestamp 1711041810
transform 0 1 21906 -1 0 22718
box -296 -734 296 766
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XMp_bias
timestamp 1711036998
transform 0 1 21873 -1 0 19854
box -296 -1219 296 1219
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_1
timestamp 1711037431
transform 0 1 21914 1 0 20509
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_2
timestamp 1711037431
transform 0 1 21914 1 0 21017
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_3
timestamp 1711037431
transform 0 1 21914 1 0 21525
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bias_4
timestamp 1711037431
transform 0 1 21914 1 0 22033
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_bot
timestamp 1711037431
transform 0 1 21914 -1 0 18185
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_mid
timestamp 1711037431
transform 0 1 21914 -1 0 18693
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_5KDBRF  XR_top
timestamp 1711037431
transform 0 1 21914 -1 0 19201
box -307 -1282 307 1282
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 DO_OUT
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 V_DISCH_O
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 V_THRESH_I
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 V_TRIG_B_I
port 5 nsew
<< end >>
