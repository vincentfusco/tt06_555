magic
tech sky130A
magscale 1 2
timestamp 1710860902
<< error_p >>
rect -77 1199 -19 1205
rect -77 1165 -65 1199
rect -77 1159 -19 1165
rect 19 71 77 77
rect 19 37 31 71
rect 19 31 77 37
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 19 -77 77 -71
rect -77 -1165 -19 -1159
rect -77 -1199 -65 -1165
rect -77 -1205 -19 -1199
<< nwell >>
rect -263 -1337 263 1337
<< pmos >>
rect -63 118 -33 1118
rect 33 118 63 1118
rect -63 -1118 -33 -118
rect 33 -1118 63 -118
<< pdiff >>
rect -125 1106 -63 1118
rect -125 130 -113 1106
rect -79 130 -63 1106
rect -125 118 -63 130
rect -33 1106 33 1118
rect -33 130 -17 1106
rect 17 130 33 1106
rect -33 118 33 130
rect 63 1106 125 1118
rect 63 130 79 1106
rect 113 130 125 1106
rect 63 118 125 130
rect -125 -130 -63 -118
rect -125 -1106 -113 -130
rect -79 -1106 -63 -130
rect -125 -1118 -63 -1106
rect -33 -130 33 -118
rect -33 -1106 -17 -130
rect 17 -1106 33 -130
rect -33 -1118 33 -1106
rect 63 -130 125 -118
rect 63 -1106 79 -130
rect 113 -1106 125 -130
rect 63 -1118 125 -1106
<< pdiffc >>
rect -113 130 -79 1106
rect -17 130 17 1106
rect 79 130 113 1106
rect -113 -1106 -79 -130
rect -17 -1106 17 -130
rect 79 -1106 113 -130
<< nsubdiff >>
rect -227 1267 -131 1301
rect 131 1267 227 1301
rect -227 1205 -193 1267
rect 193 1205 227 1267
rect -227 -1267 -193 -1205
rect 193 -1267 227 -1205
rect -227 -1301 -131 -1267
rect 131 -1301 227 -1267
<< nsubdiffcont >>
rect -131 1267 131 1301
rect -227 -1205 -193 1205
rect 193 -1205 227 1205
rect -131 -1301 131 -1267
<< poly >>
rect -81 1199 -15 1215
rect -81 1165 -65 1199
rect -31 1165 -15 1199
rect -81 1149 -15 1165
rect -63 1118 -33 1149
rect 33 1118 63 1144
rect -63 92 -33 118
rect 33 87 63 118
rect 15 71 81 87
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 15 -87 81 -71
rect -63 -118 -33 -92
rect 33 -118 63 -87
rect -63 -1149 -33 -1118
rect 33 -1144 63 -1118
rect -81 -1165 -15 -1149
rect -81 -1199 -65 -1165
rect -31 -1199 -15 -1165
rect -81 -1215 -15 -1199
<< polycont >>
rect -65 1165 -31 1199
rect 31 37 65 71
rect 31 -71 65 -37
rect -65 -1199 -31 -1165
<< locali >>
rect -227 1267 -131 1301
rect 131 1267 227 1301
rect -227 1205 -193 1267
rect 193 1205 227 1267
rect -81 1165 -65 1199
rect -31 1165 -15 1199
rect -113 1106 -79 1122
rect -113 114 -79 130
rect -17 1106 17 1122
rect -17 114 17 130
rect 79 1106 113 1122
rect 79 114 113 130
rect 15 37 31 71
rect 65 37 81 71
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -113 -130 -79 -114
rect -113 -1122 -79 -1106
rect -17 -130 17 -114
rect -17 -1122 17 -1106
rect 79 -130 113 -114
rect 79 -1122 113 -1106
rect -81 -1199 -65 -1165
rect -31 -1199 -15 -1165
rect -227 -1267 -193 -1205
rect 193 -1267 227 -1205
rect -227 -1301 -131 -1267
rect 131 -1301 227 -1267
<< viali >>
rect -65 1165 -31 1199
rect -113 130 -79 1106
rect -17 130 17 1106
rect 79 130 113 1106
rect 31 37 65 71
rect 31 -71 65 -37
rect -113 -1106 -79 -130
rect -17 -1106 17 -130
rect 79 -1106 113 -130
rect -65 -1199 -31 -1165
<< metal1 >>
rect -77 1199 -19 1205
rect -77 1165 -65 1199
rect -31 1165 -19 1199
rect -77 1159 -19 1165
rect -119 1106 -73 1118
rect -119 130 -113 1106
rect -79 130 -73 1106
rect -119 118 -73 130
rect -23 1106 23 1118
rect -23 130 -17 1106
rect 17 130 23 1106
rect -23 118 23 130
rect 73 1106 119 1118
rect 73 130 79 1106
rect 113 130 119 1106
rect 73 118 119 130
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect -119 -130 -73 -118
rect -119 -1106 -113 -130
rect -79 -1106 -73 -130
rect -119 -1118 -73 -1106
rect -23 -130 23 -118
rect -23 -1106 -17 -130
rect 17 -1106 23 -130
rect -23 -1118 23 -1106
rect 73 -130 119 -118
rect 73 -1106 79 -130
rect 113 -1106 119 -130
rect 73 -1118 119 -1106
rect -77 -1165 -19 -1159
rect -77 -1199 -65 -1165
rect -31 -1199 -19 -1165
rect -77 -1205 -19 -1199
<< properties >>
string FIXED_BBOX -210 -1284 210 1284
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
