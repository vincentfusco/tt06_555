magic
tech sky130A
magscale 1 2
timestamp 1710979170
<< error_p >>
rect -29 1775 29 1781
rect -29 1741 -17 1775
rect -29 1735 29 1741
rect -29 1581 29 1587
rect -29 1547 -17 1581
rect -29 1541 29 1547
rect -29 1473 29 1479
rect -29 1439 -17 1473
rect -29 1433 29 1439
rect -29 1279 29 1285
rect -29 1245 -17 1279
rect -29 1239 29 1245
rect -29 1171 29 1177
rect -29 1137 -17 1171
rect -29 1131 29 1137
rect -29 977 29 983
rect -29 943 -17 977
rect -29 937 29 943
rect -29 869 29 875
rect -29 835 -17 869
rect -29 829 29 835
rect -29 675 29 681
rect -29 641 -17 675
rect -29 635 29 641
rect -29 567 29 573
rect -29 533 -17 567
rect -29 527 29 533
rect -29 373 29 379
rect -29 339 -17 373
rect -29 333 29 339
rect -29 265 29 271
rect -29 231 -17 265
rect -29 225 29 231
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -231 29 -225
rect -29 -265 -17 -231
rect -29 -271 29 -265
rect -29 -339 29 -333
rect -29 -373 -17 -339
rect -29 -379 29 -373
rect -29 -533 29 -527
rect -29 -567 -17 -533
rect -29 -573 29 -567
rect -29 -641 29 -635
rect -29 -675 -17 -641
rect -29 -681 29 -675
rect -29 -835 29 -829
rect -29 -869 -17 -835
rect -29 -875 29 -869
rect -29 -943 29 -937
rect -29 -977 -17 -943
rect -29 -983 29 -977
rect -29 -1137 29 -1131
rect -29 -1171 -17 -1137
rect -29 -1177 29 -1171
rect -29 -1245 29 -1239
rect -29 -1279 -17 -1245
rect -29 -1285 29 -1279
rect -29 -1439 29 -1433
rect -29 -1473 -17 -1439
rect -29 -1479 29 -1473
rect -29 -1547 29 -1541
rect -29 -1581 -17 -1547
rect -29 -1587 29 -1581
rect -29 -1741 29 -1735
rect -29 -1775 -17 -1741
rect -29 -1781 29 -1775
<< pwell >>
rect -211 -1913 211 1913
<< nmos >>
rect -15 1619 15 1703
rect -15 1317 15 1401
rect -15 1015 15 1099
rect -15 713 15 797
rect -15 411 15 495
rect -15 109 15 193
rect -15 -193 15 -109
rect -15 -495 15 -411
rect -15 -797 15 -713
rect -15 -1099 15 -1015
rect -15 -1401 15 -1317
rect -15 -1703 15 -1619
<< ndiff >>
rect -73 1691 -15 1703
rect -73 1631 -61 1691
rect -27 1631 -15 1691
rect -73 1619 -15 1631
rect 15 1691 73 1703
rect 15 1631 27 1691
rect 61 1631 73 1691
rect 15 1619 73 1631
rect -73 1389 -15 1401
rect -73 1329 -61 1389
rect -27 1329 -15 1389
rect -73 1317 -15 1329
rect 15 1389 73 1401
rect 15 1329 27 1389
rect 61 1329 73 1389
rect 15 1317 73 1329
rect -73 1087 -15 1099
rect -73 1027 -61 1087
rect -27 1027 -15 1087
rect -73 1015 -15 1027
rect 15 1087 73 1099
rect 15 1027 27 1087
rect 61 1027 73 1087
rect 15 1015 73 1027
rect -73 785 -15 797
rect -73 725 -61 785
rect -27 725 -15 785
rect -73 713 -15 725
rect 15 785 73 797
rect 15 725 27 785
rect 61 725 73 785
rect 15 713 73 725
rect -73 483 -15 495
rect -73 423 -61 483
rect -27 423 -15 483
rect -73 411 -15 423
rect 15 483 73 495
rect 15 423 27 483
rect 61 423 73 483
rect 15 411 73 423
rect -73 181 -15 193
rect -73 121 -61 181
rect -27 121 -15 181
rect -73 109 -15 121
rect 15 181 73 193
rect 15 121 27 181
rect 61 121 73 181
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -181 -61 -121
rect -27 -181 -15 -121
rect -73 -193 -15 -181
rect 15 -121 73 -109
rect 15 -181 27 -121
rect 61 -181 73 -121
rect 15 -193 73 -181
rect -73 -423 -15 -411
rect -73 -483 -61 -423
rect -27 -483 -15 -423
rect -73 -495 -15 -483
rect 15 -423 73 -411
rect 15 -483 27 -423
rect 61 -483 73 -423
rect 15 -495 73 -483
rect -73 -725 -15 -713
rect -73 -785 -61 -725
rect -27 -785 -15 -725
rect -73 -797 -15 -785
rect 15 -725 73 -713
rect 15 -785 27 -725
rect 61 -785 73 -725
rect 15 -797 73 -785
rect -73 -1027 -15 -1015
rect -73 -1087 -61 -1027
rect -27 -1087 -15 -1027
rect -73 -1099 -15 -1087
rect 15 -1027 73 -1015
rect 15 -1087 27 -1027
rect 61 -1087 73 -1027
rect 15 -1099 73 -1087
rect -73 -1329 -15 -1317
rect -73 -1389 -61 -1329
rect -27 -1389 -15 -1329
rect -73 -1401 -15 -1389
rect 15 -1329 73 -1317
rect 15 -1389 27 -1329
rect 61 -1389 73 -1329
rect 15 -1401 73 -1389
rect -73 -1631 -15 -1619
rect -73 -1691 -61 -1631
rect -27 -1691 -15 -1631
rect -73 -1703 -15 -1691
rect 15 -1631 73 -1619
rect 15 -1691 27 -1631
rect 61 -1691 73 -1631
rect 15 -1703 73 -1691
<< ndiffc >>
rect -61 1631 -27 1691
rect 27 1631 61 1691
rect -61 1329 -27 1389
rect 27 1329 61 1389
rect -61 1027 -27 1087
rect 27 1027 61 1087
rect -61 725 -27 785
rect 27 725 61 785
rect -61 423 -27 483
rect 27 423 61 483
rect -61 121 -27 181
rect 27 121 61 181
rect -61 -181 -27 -121
rect 27 -181 61 -121
rect -61 -483 -27 -423
rect 27 -483 61 -423
rect -61 -785 -27 -725
rect 27 -785 61 -725
rect -61 -1087 -27 -1027
rect 27 -1087 61 -1027
rect -61 -1389 -27 -1329
rect 27 -1389 61 -1329
rect -61 -1691 -27 -1631
rect 27 -1691 61 -1631
<< psubdiff >>
rect -175 1843 -79 1877
rect 79 1843 175 1877
rect -175 1781 -141 1843
rect 141 1781 175 1843
rect -175 -1843 -141 -1781
rect 141 -1843 175 -1781
rect -175 -1877 -79 -1843
rect 79 -1877 175 -1843
<< psubdiffcont >>
rect -79 1843 79 1877
rect -175 -1781 -141 1781
rect 141 -1781 175 1781
rect -79 -1877 79 -1843
<< poly >>
rect -33 1775 33 1791
rect -33 1741 -17 1775
rect 17 1741 33 1775
rect -33 1725 33 1741
rect -15 1703 15 1725
rect -15 1597 15 1619
rect -33 1581 33 1597
rect -33 1547 -17 1581
rect 17 1547 33 1581
rect -33 1531 33 1547
rect -33 1473 33 1489
rect -33 1439 -17 1473
rect 17 1439 33 1473
rect -33 1423 33 1439
rect -15 1401 15 1423
rect -15 1295 15 1317
rect -33 1279 33 1295
rect -33 1245 -17 1279
rect 17 1245 33 1279
rect -33 1229 33 1245
rect -33 1171 33 1187
rect -33 1137 -17 1171
rect 17 1137 33 1171
rect -33 1121 33 1137
rect -15 1099 15 1121
rect -15 993 15 1015
rect -33 977 33 993
rect -33 943 -17 977
rect 17 943 33 977
rect -33 927 33 943
rect -33 869 33 885
rect -33 835 -17 869
rect 17 835 33 869
rect -33 819 33 835
rect -15 797 15 819
rect -15 691 15 713
rect -33 675 33 691
rect -33 641 -17 675
rect 17 641 33 675
rect -33 625 33 641
rect -33 567 33 583
rect -33 533 -17 567
rect 17 533 33 567
rect -33 517 33 533
rect -15 495 15 517
rect -15 389 15 411
rect -33 373 33 389
rect -33 339 -17 373
rect 17 339 33 373
rect -33 323 33 339
rect -33 265 33 281
rect -33 231 -17 265
rect 17 231 33 265
rect -33 215 33 231
rect -15 193 15 215
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -215 15 -193
rect -33 -231 33 -215
rect -33 -265 -17 -231
rect 17 -265 33 -231
rect -33 -281 33 -265
rect -33 -339 33 -323
rect -33 -373 -17 -339
rect 17 -373 33 -339
rect -33 -389 33 -373
rect -15 -411 15 -389
rect -15 -517 15 -495
rect -33 -533 33 -517
rect -33 -567 -17 -533
rect 17 -567 33 -533
rect -33 -583 33 -567
rect -33 -641 33 -625
rect -33 -675 -17 -641
rect 17 -675 33 -641
rect -33 -691 33 -675
rect -15 -713 15 -691
rect -15 -819 15 -797
rect -33 -835 33 -819
rect -33 -869 -17 -835
rect 17 -869 33 -835
rect -33 -885 33 -869
rect -33 -943 33 -927
rect -33 -977 -17 -943
rect 17 -977 33 -943
rect -33 -993 33 -977
rect -15 -1015 15 -993
rect -15 -1121 15 -1099
rect -33 -1137 33 -1121
rect -33 -1171 -17 -1137
rect 17 -1171 33 -1137
rect -33 -1187 33 -1171
rect -33 -1245 33 -1229
rect -33 -1279 -17 -1245
rect 17 -1279 33 -1245
rect -33 -1295 33 -1279
rect -15 -1317 15 -1295
rect -15 -1423 15 -1401
rect -33 -1439 33 -1423
rect -33 -1473 -17 -1439
rect 17 -1473 33 -1439
rect -33 -1489 33 -1473
rect -33 -1547 33 -1531
rect -33 -1581 -17 -1547
rect 17 -1581 33 -1547
rect -33 -1597 33 -1581
rect -15 -1619 15 -1597
rect -15 -1725 15 -1703
rect -33 -1741 33 -1725
rect -33 -1775 -17 -1741
rect 17 -1775 33 -1741
rect -33 -1791 33 -1775
<< polycont >>
rect -17 1741 17 1775
rect -17 1547 17 1581
rect -17 1439 17 1473
rect -17 1245 17 1279
rect -17 1137 17 1171
rect -17 943 17 977
rect -17 835 17 869
rect -17 641 17 675
rect -17 533 17 567
rect -17 339 17 373
rect -17 231 17 265
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -265 17 -231
rect -17 -373 17 -339
rect -17 -567 17 -533
rect -17 -675 17 -641
rect -17 -869 17 -835
rect -17 -977 17 -943
rect -17 -1171 17 -1137
rect -17 -1279 17 -1245
rect -17 -1473 17 -1439
rect -17 -1581 17 -1547
rect -17 -1775 17 -1741
<< locali >>
rect -175 1843 -79 1877
rect 79 1843 175 1877
rect -175 1781 -141 1843
rect 141 1781 175 1843
rect -33 1741 -17 1775
rect 17 1741 33 1775
rect -61 1691 -27 1707
rect -61 1615 -27 1631
rect 27 1691 61 1707
rect 27 1615 61 1631
rect -33 1547 -17 1581
rect 17 1547 33 1581
rect -33 1439 -17 1473
rect 17 1439 33 1473
rect -61 1389 -27 1405
rect -61 1313 -27 1329
rect 27 1389 61 1405
rect 27 1313 61 1329
rect -33 1245 -17 1279
rect 17 1245 33 1279
rect -33 1137 -17 1171
rect 17 1137 33 1171
rect -61 1087 -27 1103
rect -61 1011 -27 1027
rect 27 1087 61 1103
rect 27 1011 61 1027
rect -33 943 -17 977
rect 17 943 33 977
rect -33 835 -17 869
rect 17 835 33 869
rect -61 785 -27 801
rect -61 709 -27 725
rect 27 785 61 801
rect 27 709 61 725
rect -33 641 -17 675
rect 17 641 33 675
rect -33 533 -17 567
rect 17 533 33 567
rect -61 483 -27 499
rect -61 407 -27 423
rect 27 483 61 499
rect 27 407 61 423
rect -33 339 -17 373
rect 17 339 33 373
rect -33 231 -17 265
rect 17 231 33 265
rect -61 181 -27 197
rect -61 105 -27 121
rect 27 181 61 197
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -197 -27 -181
rect 27 -121 61 -105
rect 27 -197 61 -181
rect -33 -265 -17 -231
rect 17 -265 33 -231
rect -33 -373 -17 -339
rect 17 -373 33 -339
rect -61 -423 -27 -407
rect -61 -499 -27 -483
rect 27 -423 61 -407
rect 27 -499 61 -483
rect -33 -567 -17 -533
rect 17 -567 33 -533
rect -33 -675 -17 -641
rect 17 -675 33 -641
rect -61 -725 -27 -709
rect -61 -801 -27 -785
rect 27 -725 61 -709
rect 27 -801 61 -785
rect -33 -869 -17 -835
rect 17 -869 33 -835
rect -33 -977 -17 -943
rect 17 -977 33 -943
rect -61 -1027 -27 -1011
rect -61 -1103 -27 -1087
rect 27 -1027 61 -1011
rect 27 -1103 61 -1087
rect -33 -1171 -17 -1137
rect 17 -1171 33 -1137
rect -33 -1279 -17 -1245
rect 17 -1279 33 -1245
rect -61 -1329 -27 -1313
rect -61 -1405 -27 -1389
rect 27 -1329 61 -1313
rect 27 -1405 61 -1389
rect -33 -1473 -17 -1439
rect 17 -1473 33 -1439
rect -33 -1581 -17 -1547
rect 17 -1581 33 -1547
rect -61 -1631 -27 -1615
rect -61 -1707 -27 -1691
rect 27 -1631 61 -1615
rect 27 -1707 61 -1691
rect -33 -1775 -17 -1741
rect 17 -1775 33 -1741
rect -175 -1843 -141 -1781
rect 141 -1843 175 -1781
rect -175 -1877 -79 -1843
rect 79 -1877 175 -1843
<< viali >>
rect -17 1741 17 1775
rect -61 1631 -27 1691
rect 27 1631 61 1691
rect -17 1547 17 1581
rect -17 1439 17 1473
rect -61 1329 -27 1389
rect 27 1329 61 1389
rect -17 1245 17 1279
rect -17 1137 17 1171
rect -61 1027 -27 1087
rect 27 1027 61 1087
rect -17 943 17 977
rect -17 835 17 869
rect -61 725 -27 785
rect 27 725 61 785
rect -17 641 17 675
rect -17 533 17 567
rect -61 423 -27 483
rect 27 423 61 483
rect -17 339 17 373
rect -17 231 17 265
rect -61 121 -27 181
rect 27 121 61 181
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -181 -27 -121
rect 27 -181 61 -121
rect -17 -265 17 -231
rect -17 -373 17 -339
rect -61 -483 -27 -423
rect 27 -483 61 -423
rect -17 -567 17 -533
rect -17 -675 17 -641
rect -61 -785 -27 -725
rect 27 -785 61 -725
rect -17 -869 17 -835
rect -17 -977 17 -943
rect -61 -1087 -27 -1027
rect 27 -1087 61 -1027
rect -17 -1171 17 -1137
rect -17 -1279 17 -1245
rect -61 -1389 -27 -1329
rect 27 -1389 61 -1329
rect -17 -1473 17 -1439
rect -17 -1581 17 -1547
rect -61 -1691 -27 -1631
rect 27 -1691 61 -1631
rect -17 -1775 17 -1741
<< metal1 >>
rect -29 1775 29 1781
rect -29 1741 -17 1775
rect 17 1741 29 1775
rect -29 1735 29 1741
rect -67 1691 -21 1703
rect -67 1631 -61 1691
rect -27 1631 -21 1691
rect -67 1619 -21 1631
rect 21 1691 67 1703
rect 21 1631 27 1691
rect 61 1631 67 1691
rect 21 1619 67 1631
rect -29 1581 29 1587
rect -29 1547 -17 1581
rect 17 1547 29 1581
rect -29 1541 29 1547
rect -29 1473 29 1479
rect -29 1439 -17 1473
rect 17 1439 29 1473
rect -29 1433 29 1439
rect -67 1389 -21 1401
rect -67 1329 -61 1389
rect -27 1329 -21 1389
rect -67 1317 -21 1329
rect 21 1389 67 1401
rect 21 1329 27 1389
rect 61 1329 67 1389
rect 21 1317 67 1329
rect -29 1279 29 1285
rect -29 1245 -17 1279
rect 17 1245 29 1279
rect -29 1239 29 1245
rect -29 1171 29 1177
rect -29 1137 -17 1171
rect 17 1137 29 1171
rect -29 1131 29 1137
rect -67 1087 -21 1099
rect -67 1027 -61 1087
rect -27 1027 -21 1087
rect -67 1015 -21 1027
rect 21 1087 67 1099
rect 21 1027 27 1087
rect 61 1027 67 1087
rect 21 1015 67 1027
rect -29 977 29 983
rect -29 943 -17 977
rect 17 943 29 977
rect -29 937 29 943
rect -29 869 29 875
rect -29 835 -17 869
rect 17 835 29 869
rect -29 829 29 835
rect -67 785 -21 797
rect -67 725 -61 785
rect -27 725 -21 785
rect -67 713 -21 725
rect 21 785 67 797
rect 21 725 27 785
rect 61 725 67 785
rect 21 713 67 725
rect -29 675 29 681
rect -29 641 -17 675
rect 17 641 29 675
rect -29 635 29 641
rect -29 567 29 573
rect -29 533 -17 567
rect 17 533 29 567
rect -29 527 29 533
rect -67 483 -21 495
rect -67 423 -61 483
rect -27 423 -21 483
rect -67 411 -21 423
rect 21 483 67 495
rect 21 423 27 483
rect 61 423 67 483
rect 21 411 67 423
rect -29 373 29 379
rect -29 339 -17 373
rect 17 339 29 373
rect -29 333 29 339
rect -29 265 29 271
rect -29 231 -17 265
rect 17 231 29 265
rect -29 225 29 231
rect -67 181 -21 193
rect -67 121 -61 181
rect -27 121 -21 181
rect -67 109 -21 121
rect 21 181 67 193
rect 21 121 27 181
rect 61 121 67 181
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -181 -61 -121
rect -27 -181 -21 -121
rect -67 -193 -21 -181
rect 21 -121 67 -109
rect 21 -181 27 -121
rect 61 -181 67 -121
rect 21 -193 67 -181
rect -29 -231 29 -225
rect -29 -265 -17 -231
rect 17 -265 29 -231
rect -29 -271 29 -265
rect -29 -339 29 -333
rect -29 -373 -17 -339
rect 17 -373 29 -339
rect -29 -379 29 -373
rect -67 -423 -21 -411
rect -67 -483 -61 -423
rect -27 -483 -21 -423
rect -67 -495 -21 -483
rect 21 -423 67 -411
rect 21 -483 27 -423
rect 61 -483 67 -423
rect 21 -495 67 -483
rect -29 -533 29 -527
rect -29 -567 -17 -533
rect 17 -567 29 -533
rect -29 -573 29 -567
rect -29 -641 29 -635
rect -29 -675 -17 -641
rect 17 -675 29 -641
rect -29 -681 29 -675
rect -67 -725 -21 -713
rect -67 -785 -61 -725
rect -27 -785 -21 -725
rect -67 -797 -21 -785
rect 21 -725 67 -713
rect 21 -785 27 -725
rect 61 -785 67 -725
rect 21 -797 67 -785
rect -29 -835 29 -829
rect -29 -869 -17 -835
rect 17 -869 29 -835
rect -29 -875 29 -869
rect -29 -943 29 -937
rect -29 -977 -17 -943
rect 17 -977 29 -943
rect -29 -983 29 -977
rect -67 -1027 -21 -1015
rect -67 -1087 -61 -1027
rect -27 -1087 -21 -1027
rect -67 -1099 -21 -1087
rect 21 -1027 67 -1015
rect 21 -1087 27 -1027
rect 61 -1087 67 -1027
rect 21 -1099 67 -1087
rect -29 -1137 29 -1131
rect -29 -1171 -17 -1137
rect 17 -1171 29 -1137
rect -29 -1177 29 -1171
rect -29 -1245 29 -1239
rect -29 -1279 -17 -1245
rect 17 -1279 29 -1245
rect -29 -1285 29 -1279
rect -67 -1329 -21 -1317
rect -67 -1389 -61 -1329
rect -27 -1389 -21 -1329
rect -67 -1401 -21 -1389
rect 21 -1329 67 -1317
rect 21 -1389 27 -1329
rect 61 -1389 67 -1329
rect 21 -1401 67 -1389
rect -29 -1439 29 -1433
rect -29 -1473 -17 -1439
rect 17 -1473 29 -1439
rect -29 -1479 29 -1473
rect -29 -1547 29 -1541
rect -29 -1581 -17 -1547
rect 17 -1581 29 -1547
rect -29 -1587 29 -1581
rect -67 -1631 -21 -1619
rect -67 -1691 -61 -1631
rect -27 -1691 -21 -1631
rect -67 -1703 -21 -1691
rect 21 -1631 67 -1619
rect 21 -1691 27 -1631
rect 61 -1691 67 -1631
rect 21 -1703 67 -1691
rect -29 -1741 29 -1735
rect -29 -1775 -17 -1741
rect 17 -1775 29 -1741
rect -29 -1781 29 -1775
<< properties >>
string FIXED_BBOX -158 -1860 158 1860
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 12 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
