* SPICE3 file created from tt_um_vaf_555_timer.ext - technology: sky130A

.subckt tt_um_vaf_555_timer clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VPWR VGND
C0 ua[1] VPWR 3.561736f
C1 VPWR X_TIMER/X_COMP_P_BOTTOM/out_left 6.370519f
C2 ua[0] X_TIMER/X_COMP_P_TOP/tail 2.920444f
C3 ui_in[0] X_TIMER/X_SR_LATCH/IN_R 3.252836f
C4 X_TIMER/X_COMP_P_TOP/tail X_TIMER/X_COMP_P_TOP/latch_left 8.829929f
C5 X_TIMER/X_COMP_P_BOTTOM/latch_left X_TIMER/X_COMP_P_BOTTOM/tail 8.827988f
C6 VPWR X_TIMER/X_SR_LATCH/IN_S 3.474115f
C7 X_TIMER/v1p2 X_TIMER/X_COMP_P_TOP/latch_right 3.535094f
C8 uo_out[0] VPWR 8.463964f
C9 VPWR X_TIMER/bias_p 12.319203f
C10 X_TIMER/X_COMP_P_BOTTOM/latch_left X_TIMER/X_COMP_P_BOTTOM/latch_right 5.38251f
C11 X_TIMER/X_COMP_P_BOTTOM/tail X_TIMER/X_COMP_P_BOTTOM/latch_right 8.893079f
C12 X_TIMER/X_COMP_P_TOP/tail X_TIMER/X_COMP_P_TOP/latch_right 8.894202f
C13 ua[0] ua[1] 10.74292f
C14 ua[1] X_TIMER/X_COMP_P_BOTTOM/latch_right 3.575976f
C15 ua[1] ua[2] 4.93575f
C16 X_TIMER/X_COMP_P_TOP/latch_left X_TIMER/X_COMP_P_TOP/latch_right 5.38251f
C17 VPWR X_TIMER/v0p6 5.940137f
C18 VPWR X_TIMER/X_SR_LATCH/IN_R 4.52376f
C19 X_TIMER/v0p6 X_TIMER/X_COMP_P_BOTTOM/tail 2.674759f
C20 uo_out[0] ui_in[0] 19.735884f
C21 X_TIMER/v1p2 VPWR 3.828327f
C22 X_TIMER/X_COMP_P_TOP/tail VPWR 5.099898f
C23 VPWR X_TIMER/X_COMP_P_BOTTOM/tail 5.617589f
C24 ua[0] VPWR 5.198981f
C25 X_TIMER/X_COMP_P_TOP/out_left VPWR 6.353149f
XX_TIMER ua[0] ua[1] ui_in[0] uo_out[0] ua[2] VPWR VGND timer_core
C26 X_TIMER/v1p2 VGND 3.173445f
C27 X_TIMER/v0p6 VGND 2.301639f
C28 X_TIMER/bias_n VGND 2.762814f **FLOATING
C29 uo_out[0] VGND 10.320412f
C30 ua[2] VGND 17.301718f
C31 X_TIMER/out_inv3 VGND 4.323294f
C32 ua[0] VGND 17.07561f
C33 X_TIMER/X_COMP_P_TOP/latch_right VGND 6.317735f
C34 X_TIMER/X_COMP_P_TOP/out_left VGND 3.664091f
C35 X_TIMER/X_COMP_P_TOP/latch_left VGND 6.153733f
C36 ua[1] VGND 12.375967f
C37 X_TIMER/bias_p VGND 2.868942f
C38 X_TIMER/X_COMP_P_BOTTOM/latch_right VGND 6.412793f
C39 X_TIMER/X_COMP_P_BOTTOM/out_left VGND 3.668321f
C40 X_TIMER/X_COMP_P_BOTTOM/latch_left VGND 6.207313f
C41 ui_in[0] VGND 18.061064f
C42 VPWR VGND 0.113984p
C43 X_TIMER/X_SR_LATCH/IN_S VGND 10.724534f
C44 X_TIMER/X_SR_LATCH/IN_R VGND 13.356827f
.ends
